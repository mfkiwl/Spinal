// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : Plic
// Git hash  : adf552d8f500e7419fff395b7049228e4bc5de26



module Plic (
  input      [23:0]   io_apb_PADDR,
  input      [0:0]    io_apb_PSEL,
  input               io_apb_PENABLE,
  output reg          io_apb_PREADY,
  input               io_apb_PWRITE,
  input      [31:0]   io_apb_PWDATA,
  output reg [31:0]   io_apb_PRDATA,
  output              io_apb_PSLVERROR,
  input      [34:0]   io_sources,
  output     [2:0]    io_targets,
  input               clk,
  input               reset
);
  wire                _zz_708;
  wire       [0:0]    _zz_709;
  wire       [0:0]    _zz_710;
  wire       [0:0]    _zz_711;
  wire       [0:0]    _zz_712;
  wire       [0:0]    _zz_713;
  wire       [0:0]    _zz_714;
  wire       [0:0]    _zz_715;
  wire       [0:0]    _zz_716;
  wire       [0:0]    _zz_717;
  wire       [0:0]    _zz_718;
  wire       [0:0]    _zz_719;
  wire       [0:0]    _zz_720;
  wire       [0:0]    _zz_721;
  wire       [0:0]    _zz_722;
  wire       [0:0]    _zz_723;
  wire       [0:0]    _zz_724;
  wire       [0:0]    _zz_725;
  wire       [0:0]    _zz_726;
  wire       [0:0]    _zz_727;
  wire       [0:0]    _zz_728;
  wire       [0:0]    _zz_729;
  wire       [0:0]    _zz_730;
  wire       [0:0]    _zz_731;
  wire       [0:0]    _zz_732;
  wire       [0:0]    _zz_733;
  wire       [0:0]    _zz_734;
  wire       [0:0]    _zz_735;
  wire       [0:0]    _zz_736;
  wire       [0:0]    _zz_737;
  wire       [0:0]    _zz_738;
  wire       [0:0]    _zz_739;
  wire       [0:0]    _zz_740;
  wire       [0:0]    _zz_741;
  wire       [0:0]    _zz_742;
  wire       [0:0]    _zz_743;
  wire       [0:0]    _zz_744;
  wire       [0:0]    _zz_745;
  wire       [0:0]    _zz_746;
  wire       [0:0]    _zz_747;
  wire       [0:0]    _zz_748;
  wire       [0:0]    _zz_749;
  wire       [0:0]    _zz_750;
  wire       [0:0]    _zz_751;
  wire       [0:0]    _zz_752;
  wire       [0:0]    _zz_753;
  wire       [0:0]    _zz_754;
  wire       [0:0]    _zz_755;
  wire       [0:0]    _zz_756;
  wire       [0:0]    _zz_757;
  wire       [0:0]    _zz_758;
  wire       [0:0]    _zz_759;
  wire       [0:0]    _zz_760;
  wire       [0:0]    _zz_761;
  wire       [0:0]    _zz_762;
  wire       [0:0]    _zz_763;
  wire       [0:0]    _zz_764;
  wire       [0:0]    _zz_765;
  wire       [0:0]    _zz_766;
  wire       [0:0]    _zz_767;
  wire       [0:0]    _zz_768;
  wire       [0:0]    _zz_769;
  wire       [0:0]    _zz_770;
  wire       [0:0]    _zz_771;
  wire       [0:0]    _zz_772;
  wire       [0:0]    _zz_773;
  wire       [0:0]    _zz_774;
  wire       [0:0]    _zz_775;
  wire       [0:0]    _zz_776;
  wire       [0:0]    _zz_777;
  wire       [0:0]    _zz_778;
  wire       [0:0]    _zz_779;
  wire       [0:0]    _zz_780;
  wire       [0:0]    _zz_781;
  wire       [0:0]    _zz_782;
  wire       [0:0]    _zz_783;
  wire       [0:0]    _zz_784;
  wire       [0:0]    _zz_785;
  wire       [0:0]    _zz_786;
  wire       [0:0]    _zz_787;
  wire       [0:0]    _zz_788;
  wire       [0:0]    _zz_789;
  wire       [0:0]    _zz_790;
  wire       [0:0]    _zz_791;
  wire       [0:0]    _zz_792;
  wire       [0:0]    _zz_793;
  wire       [0:0]    _zz_794;
  wire       [0:0]    _zz_795;
  wire       [0:0]    _zz_796;
  wire       [0:0]    _zz_797;
  wire       [0:0]    _zz_798;
  wire       [0:0]    _zz_799;
  wire       [0:0]    _zz_800;
  wire       [0:0]    _zz_801;
  wire       [0:0]    _zz_802;
  wire       [0:0]    _zz_803;
  wire       [0:0]    _zz_804;
  wire       [0:0]    _zz_805;
  wire       [0:0]    _zz_806;
  wire       [0:0]    _zz_807;
  wire       [0:0]    _zz_808;
  wire       [0:0]    _zz_809;
  wire       [0:0]    _zz_810;
  wire       [0:0]    _zz_811;
  wire       [0:0]    _zz_812;
  wire       [0:0]    _zz_813;
  wire       [6:0]    _zz_814;
  wire       [6:0]    _zz_815;
  wire       [6:0]    _zz_816;
  wire       [6:0]    _zz_817;
  wire       [6:0]    _zz_818;
  wire       [6:0]    _zz_819;
  wire       [6:0]    _zz_820;
  wire       [6:0]    _zz_821;
  wire       [6:0]    _zz_822;
  wire       [6:0]    _zz_823;
  wire       [6:0]    _zz_824;
  wire       [6:0]    _zz_825;
  wire       [6:0]    _zz_826;
  wire       [6:0]    _zz_827;
  wire       [6:0]    _zz_828;
  wire       [6:0]    _zz_829;
  wire       [6:0]    _zz_830;
  wire       [6:0]    _zz_831;
  wire       [6:0]    _zz_832;
  wire       [6:0]    _zz_833;
  wire       [6:0]    _zz_834;
  wire       [6:0]    _zz_835;
  wire       [6:0]    _zz_836;
  wire       [6:0]    _zz_837;
  wire       [6:0]    _zz_838;
  wire       [6:0]    _zz_839;
  wire       [6:0]    _zz_840;
  wire       [6:0]    _zz_841;
  wire       [6:0]    _zz_842;
  wire       [6:0]    _zz_843;
  wire       [6:0]    _zz_844;
  wire       [6:0]    _zz_845;
  wire       [6:0]    _zz_846;
  wire       [6:0]    _zz_847;
  wire       [6:0]    _zz_848;
  wire       [6:0]    _zz_849;
  wire       [6:0]    _zz_850;
  wire       [6:0]    _zz_851;
  wire       [6:0]    _zz_852;
  wire       [6:0]    _zz_853;
  wire       [6:0]    _zz_854;
  wire       [6:0]    _zz_855;
  wire       [6:0]    _zz_856;
  wire       [6:0]    _zz_857;
  wire       [6:0]    _zz_858;
  wire       [6:0]    _zz_859;
  wire       [6:0]    _zz_860;
  wire       [6:0]    _zz_861;
  wire       [6:0]    _zz_862;
  wire       [6:0]    _zz_863;
  wire       [6:0]    _zz_864;
  wire       [6:0]    _zz_865;
  wire       [6:0]    _zz_866;
  wire       [6:0]    _zz_867;
  wire       [6:0]    _zz_868;
  wire       [6:0]    _zz_869;
  wire       [6:0]    _zz_870;
  wire       [6:0]    _zz_871;
  wire       [6:0]    _zz_872;
  wire       [6:0]    _zz_873;
  wire       [6:0]    _zz_874;
  wire       [6:0]    _zz_875;
  wire       [6:0]    _zz_876;
  wire       [6:0]    _zz_877;
  wire       [6:0]    _zz_878;
  wire       [6:0]    _zz_879;
  wire       [6:0]    _zz_880;
  wire       [6:0]    _zz_881;
  wire       [6:0]    _zz_882;
  wire       [6:0]    _zz_883;
  wire       [6:0]    _zz_884;
  wire       [6:0]    _zz_885;
  wire       [6:0]    _zz_886;
  wire       [6:0]    _zz_887;
  wire       [6:0]    _zz_888;
  wire       [6:0]    _zz_889;
  wire       [6:0]    _zz_890;
  wire       [6:0]    _zz_891;
  wire       [6:0]    _zz_892;
  wire       [6:0]    _zz_893;
  wire       [6:0]    _zz_894;
  wire       [6:0]    _zz_895;
  wire       [6:0]    _zz_896;
  wire       [6:0]    _zz_897;
  wire       [6:0]    _zz_898;
  wire       [6:0]    _zz_899;
  wire       [6:0]    _zz_900;
  wire       [6:0]    _zz_901;
  wire                _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire       [1:0]    gateways_0_priority;
  reg                 gateways_0_ip;
  reg                 gateways_0_waitCompletion;
  wire       [1:0]    gateways_1_priority;
  reg                 gateways_1_ip;
  reg                 gateways_1_waitCompletion;
  wire       [1:0]    gateways_2_priority;
  reg                 gateways_2_ip;
  reg                 gateways_2_waitCompletion;
  wire       [1:0]    gateways_3_priority;
  reg                 gateways_3_ip;
  reg                 gateways_3_waitCompletion;
  wire       [1:0]    gateways_4_priority;
  reg                 gateways_4_ip;
  reg                 gateways_4_waitCompletion;
  wire       [1:0]    gateways_5_priority;
  reg                 gateways_5_ip;
  reg                 gateways_5_waitCompletion;
  wire       [1:0]    gateways_6_priority;
  reg                 gateways_6_ip;
  reg                 gateways_6_waitCompletion;
  wire       [1:0]    gateways_7_priority;
  reg                 gateways_7_ip;
  reg                 gateways_7_waitCompletion;
  wire       [1:0]    gateways_8_priority;
  reg                 gateways_8_ip;
  reg                 gateways_8_waitCompletion;
  wire       [1:0]    gateways_9_priority;
  reg                 gateways_9_ip;
  reg                 gateways_9_waitCompletion;
  wire       [1:0]    gateways_10_priority;
  reg                 gateways_10_ip;
  reg                 gateways_10_waitCompletion;
  wire       [1:0]    gateways_11_priority;
  reg                 gateways_11_ip;
  reg                 gateways_11_waitCompletion;
  wire       [1:0]    gateways_12_priority;
  reg                 gateways_12_ip;
  reg                 gateways_12_waitCompletion;
  wire       [1:0]    gateways_13_priority;
  reg                 gateways_13_ip;
  reg                 gateways_13_waitCompletion;
  wire       [1:0]    gateways_14_priority;
  reg                 gateways_14_ip;
  reg                 gateways_14_waitCompletion;
  wire       [1:0]    gateways_15_priority;
  reg                 gateways_15_ip;
  reg                 gateways_15_waitCompletion;
  wire       [1:0]    gateways_16_priority;
  reg                 gateways_16_ip;
  reg                 gateways_16_waitCompletion;
  wire       [1:0]    gateways_17_priority;
  reg                 gateways_17_ip;
  reg                 gateways_17_waitCompletion;
  wire       [1:0]    gateways_18_priority;
  reg                 gateways_18_ip;
  reg                 gateways_18_waitCompletion;
  wire       [1:0]    gateways_19_priority;
  reg                 gateways_19_ip;
  reg                 gateways_19_waitCompletion;
  wire       [1:0]    gateways_20_priority;
  reg                 gateways_20_ip;
  reg                 gateways_20_waitCompletion;
  wire       [1:0]    gateways_21_priority;
  reg                 gateways_21_ip;
  reg                 gateways_21_waitCompletion;
  wire       [1:0]    gateways_22_priority;
  reg                 gateways_22_ip;
  reg                 gateways_22_waitCompletion;
  wire       [1:0]    gateways_23_priority;
  reg                 gateways_23_ip;
  reg                 gateways_23_waitCompletion;
  wire       [1:0]    gateways_24_priority;
  reg                 gateways_24_ip;
  reg                 gateways_24_waitCompletion;
  wire       [1:0]    gateways_25_priority;
  reg                 gateways_25_ip;
  reg                 gateways_25_waitCompletion;
  wire       [1:0]    gateways_26_priority;
  reg                 gateways_26_ip;
  reg                 gateways_26_waitCompletion;
  wire       [1:0]    gateways_27_priority;
  reg                 gateways_27_ip;
  reg                 gateways_27_waitCompletion;
  wire       [1:0]    gateways_28_priority;
  reg                 gateways_28_ip;
  reg                 gateways_28_waitCompletion;
  wire       [1:0]    gateways_29_priority;
  reg                 gateways_29_ip;
  reg                 gateways_29_waitCompletion;
  wire       [1:0]    gateways_30_priority;
  reg                 gateways_30_ip;
  reg                 gateways_30_waitCompletion;
  wire       [1:0]    gateways_31_priority;
  reg                 gateways_31_ip;
  reg                 gateways_31_waitCompletion;
  wire       [1:0]    gateways_32_priority;
  reg                 gateways_32_ip;
  reg                 gateways_32_waitCompletion;
  wire       [1:0]    gateways_33_priority;
  reg                 gateways_33_ip;
  reg                 gateways_33_waitCompletion;
  wire       [1:0]    gateways_34_priority;
  reg                 gateways_34_ip;
  reg                 gateways_34_waitCompletion;
  wire                targets_0_ie_0;
  wire                targets_0_ie_1;
  wire                targets_0_ie_2;
  wire                targets_0_ie_3;
  wire                targets_0_ie_4;
  wire                targets_0_ie_5;
  wire                targets_0_ie_6;
  wire                targets_0_ie_7;
  wire                targets_0_ie_8;
  wire                targets_0_ie_9;
  wire                targets_0_ie_10;
  wire                targets_0_ie_11;
  wire                targets_0_ie_12;
  wire                targets_0_ie_13;
  wire                targets_0_ie_14;
  wire                targets_0_ie_15;
  wire                targets_0_ie_16;
  wire                targets_0_ie_17;
  wire                targets_0_ie_18;
  wire                targets_0_ie_19;
  wire                targets_0_ie_20;
  wire                targets_0_ie_21;
  wire                targets_0_ie_22;
  wire                targets_0_ie_23;
  wire                targets_0_ie_24;
  wire                targets_0_ie_25;
  wire                targets_0_ie_26;
  wire                targets_0_ie_27;
  wire                targets_0_ie_28;
  wire                targets_0_ie_29;
  wire                targets_0_ie_30;
  wire                targets_0_ie_31;
  wire                targets_0_ie_32;
  wire                targets_0_ie_33;
  wire                targets_0_ie_34;
  wire       [1:0]    targets_0_threshold;
  wire       [1:0]    targets_0_requests_0_priority;
  wire       [6:0]    targets_0_requests_0_id;
  wire                targets_0_requests_0_valid;
  wire       [1:0]    targets_0_requests_1_priority;
  wire       [6:0]    targets_0_requests_1_id;
  wire                targets_0_requests_1_valid;
  wire       [1:0]    targets_0_requests_2_priority;
  wire       [6:0]    targets_0_requests_2_id;
  wire                targets_0_requests_2_valid;
  wire       [1:0]    targets_0_requests_3_priority;
  wire       [6:0]    targets_0_requests_3_id;
  wire                targets_0_requests_3_valid;
  wire       [1:0]    targets_0_requests_4_priority;
  wire       [6:0]    targets_0_requests_4_id;
  wire                targets_0_requests_4_valid;
  wire       [1:0]    targets_0_requests_5_priority;
  wire       [6:0]    targets_0_requests_5_id;
  wire                targets_0_requests_5_valid;
  wire       [1:0]    targets_0_requests_6_priority;
  wire       [6:0]    targets_0_requests_6_id;
  wire                targets_0_requests_6_valid;
  wire       [1:0]    targets_0_requests_7_priority;
  wire       [6:0]    targets_0_requests_7_id;
  wire                targets_0_requests_7_valid;
  wire       [1:0]    targets_0_requests_8_priority;
  wire       [6:0]    targets_0_requests_8_id;
  wire                targets_0_requests_8_valid;
  wire       [1:0]    targets_0_requests_9_priority;
  wire       [6:0]    targets_0_requests_9_id;
  wire                targets_0_requests_9_valid;
  wire       [1:0]    targets_0_requests_10_priority;
  wire       [6:0]    targets_0_requests_10_id;
  wire                targets_0_requests_10_valid;
  wire       [1:0]    targets_0_requests_11_priority;
  wire       [6:0]    targets_0_requests_11_id;
  wire                targets_0_requests_11_valid;
  wire       [1:0]    targets_0_requests_12_priority;
  wire       [6:0]    targets_0_requests_12_id;
  wire                targets_0_requests_12_valid;
  wire       [1:0]    targets_0_requests_13_priority;
  wire       [6:0]    targets_0_requests_13_id;
  wire                targets_0_requests_13_valid;
  wire       [1:0]    targets_0_requests_14_priority;
  wire       [6:0]    targets_0_requests_14_id;
  wire                targets_0_requests_14_valid;
  wire       [1:0]    targets_0_requests_15_priority;
  wire       [6:0]    targets_0_requests_15_id;
  wire                targets_0_requests_15_valid;
  wire       [1:0]    targets_0_requests_16_priority;
  wire       [6:0]    targets_0_requests_16_id;
  wire                targets_0_requests_16_valid;
  wire       [1:0]    targets_0_requests_17_priority;
  wire       [6:0]    targets_0_requests_17_id;
  wire                targets_0_requests_17_valid;
  wire       [1:0]    targets_0_requests_18_priority;
  wire       [6:0]    targets_0_requests_18_id;
  wire                targets_0_requests_18_valid;
  wire       [1:0]    targets_0_requests_19_priority;
  wire       [6:0]    targets_0_requests_19_id;
  wire                targets_0_requests_19_valid;
  wire       [1:0]    targets_0_requests_20_priority;
  wire       [6:0]    targets_0_requests_20_id;
  wire                targets_0_requests_20_valid;
  wire       [1:0]    targets_0_requests_21_priority;
  wire       [6:0]    targets_0_requests_21_id;
  wire                targets_0_requests_21_valid;
  wire       [1:0]    targets_0_requests_22_priority;
  wire       [6:0]    targets_0_requests_22_id;
  wire                targets_0_requests_22_valid;
  wire       [1:0]    targets_0_requests_23_priority;
  wire       [6:0]    targets_0_requests_23_id;
  wire                targets_0_requests_23_valid;
  wire       [1:0]    targets_0_requests_24_priority;
  wire       [6:0]    targets_0_requests_24_id;
  wire                targets_0_requests_24_valid;
  wire       [1:0]    targets_0_requests_25_priority;
  wire       [6:0]    targets_0_requests_25_id;
  wire                targets_0_requests_25_valid;
  wire       [1:0]    targets_0_requests_26_priority;
  wire       [6:0]    targets_0_requests_26_id;
  wire                targets_0_requests_26_valid;
  wire       [1:0]    targets_0_requests_27_priority;
  wire       [6:0]    targets_0_requests_27_id;
  wire                targets_0_requests_27_valid;
  wire       [1:0]    targets_0_requests_28_priority;
  wire       [6:0]    targets_0_requests_28_id;
  wire                targets_0_requests_28_valid;
  wire       [1:0]    targets_0_requests_29_priority;
  wire       [6:0]    targets_0_requests_29_id;
  wire                targets_0_requests_29_valid;
  wire       [1:0]    targets_0_requests_30_priority;
  wire       [6:0]    targets_0_requests_30_id;
  wire                targets_0_requests_30_valid;
  wire       [1:0]    targets_0_requests_31_priority;
  wire       [6:0]    targets_0_requests_31_id;
  wire                targets_0_requests_31_valid;
  wire       [1:0]    targets_0_requests_32_priority;
  wire       [6:0]    targets_0_requests_32_id;
  wire                targets_0_requests_32_valid;
  wire       [1:0]    targets_0_requests_33_priority;
  wire       [6:0]    targets_0_requests_33_id;
  wire                targets_0_requests_33_valid;
  wire       [1:0]    targets_0_requests_34_priority;
  wire       [6:0]    targets_0_requests_34_id;
  wire                targets_0_requests_34_valid;
  wire       [1:0]    targets_0_requests_35_priority;
  wire       [6:0]    targets_0_requests_35_id;
  wire                targets_0_requests_35_valid;
  wire                _zz_36;
  wire       [1:0]    _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire       [1:0]    _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire       [1:0]    _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire       [1:0]    _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire       [1:0]    _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire       [1:0]    _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire       [1:0]    _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire       [1:0]    _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire       [1:0]    _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire       [1:0]    _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire       [1:0]    _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire       [1:0]    _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire       [1:0]    _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire       [1:0]    _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire       [1:0]    _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire       [1:0]    _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire       [1:0]    _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire       [1:0]    _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire       [1:0]    _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire       [1:0]    _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire       [1:0]    _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire       [1:0]    _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire       [1:0]    _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire       [1:0]    _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire       [1:0]    _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire       [1:0]    _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire       [1:0]    _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire       [1:0]    _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire       [1:0]    _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire       [1:0]    _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire       [1:0]    _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire       [1:0]    _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire       [1:0]    _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire       [1:0]    _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  reg        [1:0]    targets_0_bestRequest_priority;
  reg        [6:0]    targets_0_bestRequest_id;
  reg                 targets_0_bestRequest_valid;
  wire                targets_0_iep;
  wire       [6:0]    targets_0_claim;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire       [1:0]    _zz_174;
  wire       [1:0]    _zz_175;
  wire                _zz_176;
  wire       [1:0]    _zz_177;
  wire                _zz_178;
  wire       [1:0]    _zz_179;
  wire                _zz_180;
  wire       [1:0]    _zz_181;
  wire                _zz_182;
  wire       [1:0]    _zz_183;
  wire                _zz_184;
  wire       [1:0]    _zz_185;
  wire                _zz_186;
  wire       [1:0]    _zz_187;
  wire                _zz_188;
  wire       [1:0]    _zz_189;
  wire                _zz_190;
  wire       [1:0]    _zz_191;
  wire                _zz_192;
  wire       [1:0]    _zz_193;
  wire                _zz_194;
  wire       [1:0]    _zz_195;
  wire                _zz_196;
  wire       [1:0]    _zz_197;
  wire                _zz_198;
  wire       [1:0]    _zz_199;
  wire                _zz_200;
  wire       [1:0]    _zz_201;
  wire                _zz_202;
  wire       [1:0]    _zz_203;
  wire                _zz_204;
  wire       [1:0]    _zz_205;
  wire                _zz_206;
  wire       [1:0]    _zz_207;
  wire                _zz_208;
  wire       [1:0]    _zz_209;
  wire                _zz_210;
  wire       [1:0]    _zz_211;
  wire                _zz_212;
  wire       [1:0]    _zz_213;
  wire                _zz_214;
  wire       [1:0]    _zz_215;
  wire                _zz_216;
  wire       [1:0]    _zz_217;
  wire                _zz_218;
  wire       [1:0]    _zz_219;
  wire                _zz_220;
  wire       [1:0]    _zz_221;
  wire                _zz_222;
  wire       [1:0]    _zz_223;
  wire                _zz_224;
  wire       [1:0]    _zz_225;
  wire                _zz_226;
  wire       [1:0]    _zz_227;
  wire                _zz_228;
  wire       [1:0]    _zz_229;
  wire                _zz_230;
  wire       [1:0]    _zz_231;
  wire                _zz_232;
  wire       [1:0]    _zz_233;
  wire                _zz_234;
  wire       [1:0]    _zz_235;
  wire                _zz_236;
  wire       [1:0]    _zz_237;
  wire                _zz_238;
  wire       [1:0]    _zz_239;
  wire                _zz_240;
  wire       [1:0]    _zz_241;
  wire                _zz_242;
  wire       [1:0]    _zz_243;
  wire                _zz_244;
  wire       [1:0]    _zz_245;
  wire                _zz_246;
  wire                _zz_247;
  wire       [1:0]    _zz_248;
  wire                _zz_249;
  wire                _zz_250;
  wire       [1:0]    _zz_251;
  wire                _zz_252;
  wire                _zz_253;
  wire       [1:0]    _zz_254;
  wire                _zz_255;
  wire                _zz_256;
  wire       [1:0]    _zz_257;
  wire                _zz_258;
  wire                _zz_259;
  wire       [1:0]    _zz_260;
  wire                _zz_261;
  wire                _zz_262;
  wire       [1:0]    _zz_263;
  wire                _zz_264;
  wire                _zz_265;
  wire       [1:0]    _zz_266;
  wire                _zz_267;
  wire                _zz_268;
  wire       [1:0]    _zz_269;
  wire                _zz_270;
  wire                _zz_271;
  wire       [1:0]    _zz_272;
  wire                _zz_273;
  wire                _zz_274;
  wire       [1:0]    _zz_275;
  wire                _zz_276;
  wire                _zz_277;
  wire       [1:0]    _zz_278;
  wire                _zz_279;
  wire                _zz_280;
  wire       [1:0]    _zz_281;
  wire                _zz_282;
  wire                _zz_283;
  wire       [1:0]    _zz_284;
  wire                _zz_285;
  wire                _zz_286;
  wire       [1:0]    _zz_287;
  wire                _zz_288;
  wire                _zz_289;
  wire       [1:0]    _zz_290;
  wire                _zz_291;
  wire                _zz_292;
  wire       [1:0]    _zz_293;
  wire                _zz_294;
  wire                _zz_295;
  wire       [1:0]    _zz_296;
  wire                _zz_297;
  wire                _zz_298;
  wire       [1:0]    _zz_299;
  wire                _zz_300;
  wire                _zz_301;
  wire       [1:0]    _zz_302;
  wire                _zz_303;
  wire                _zz_304;
  wire       [1:0]    _zz_305;
  wire                _zz_306;
  wire                _zz_307;
  wire       [1:0]    _zz_308;
  wire                _zz_309;
  wire                _zz_310;
  wire       [1:0]    _zz_311;
  wire                _zz_312;
  wire                _zz_313;
  wire       [1:0]    _zz_314;
  wire                _zz_315;
  wire                _zz_316;
  wire       [1:0]    _zz_317;
  wire                _zz_318;
  wire                _zz_319;
  wire       [1:0]    _zz_320;
  wire                _zz_321;
  wire                _zz_322;
  wire       [1:0]    _zz_323;
  wire                _zz_324;
  wire                _zz_325;
  wire       [1:0]    _zz_326;
  wire                _zz_327;
  wire       [1:0]    _zz_328;
  wire                _zz_329;
  wire                _zz_330;
  wire       [1:0]    _zz_331;
  wire                _zz_332;
  wire                _zz_333;
  wire       [1:0]    _zz_334;
  wire                _zz_335;
  wire                _zz_336;
  wire       [1:0]    _zz_337;
  wire                _zz_338;
  wire                _zz_339;
  wire       [1:0]    _zz_340;
  wire                _zz_341;
  wire                _zz_342;
  wire       [1:0]    _zz_343;
  wire                _zz_344;
  wire                _zz_345;
  wire       [1:0]    _zz_346;
  wire                _zz_347;
  reg        [1:0]    _zz_348;
  reg        [6:0]    _zz_349;
  wire                _zz_350;
  wire       [6:0]    _zz_351;
  wire                _zz_352;
  wire                _zz_353;
  wire                _zz_354;
  wire                _zz_355;
  wire                _zz_356;
  wire                _zz_357;
  wire                _zz_358;
  wire                _zz_359;
  wire                _zz_360;
  wire                _zz_361;
  wire                _zz_362;
  wire                _zz_363;
  wire                _zz_364;
  wire                _zz_365;
  wire                _zz_366;
  wire                _zz_367;
  wire                _zz_368;
  wire                _zz_369;
  wire                _zz_370;
  wire                _zz_371;
  wire                _zz_372;
  wire                _zz_373;
  wire                _zz_374;
  wire                _zz_375;
  wire                _zz_376;
  wire                _zz_377;
  wire                _zz_378;
  wire                _zz_379;
  wire                _zz_380;
  wire                _zz_381;
  wire                _zz_382;
  wire                _zz_383;
  wire                _zz_384;
  wire                _zz_385;
  wire                _zz_386;
  wire       [1:0]    _zz_387;
  wire       [1:0]    _zz_388;
  wire                _zz_389;
  wire       [1:0]    _zz_390;
  wire                _zz_391;
  wire       [1:0]    _zz_392;
  wire                _zz_393;
  wire       [1:0]    _zz_394;
  wire                _zz_395;
  wire       [1:0]    _zz_396;
  wire                _zz_397;
  wire       [1:0]    _zz_398;
  wire                _zz_399;
  wire       [1:0]    _zz_400;
  wire                _zz_401;
  wire       [1:0]    _zz_402;
  wire                _zz_403;
  wire       [1:0]    _zz_404;
  wire                _zz_405;
  wire       [1:0]    _zz_406;
  wire                _zz_407;
  wire       [1:0]    _zz_408;
  wire                _zz_409;
  wire       [1:0]    _zz_410;
  wire                _zz_411;
  wire       [1:0]    _zz_412;
  wire                _zz_413;
  wire       [1:0]    _zz_414;
  wire                _zz_415;
  wire       [1:0]    _zz_416;
  wire                _zz_417;
  wire       [1:0]    _zz_418;
  wire                _zz_419;
  wire       [1:0]    _zz_420;
  wire                _zz_421;
  wire       [1:0]    _zz_422;
  wire                _zz_423;
  wire       [1:0]    _zz_424;
  wire                _zz_425;
  wire       [1:0]    _zz_426;
  wire                _zz_427;
  wire       [1:0]    _zz_428;
  wire                _zz_429;
  wire       [1:0]    _zz_430;
  wire                _zz_431;
  wire       [1:0]    _zz_432;
  wire                _zz_433;
  wire       [1:0]    _zz_434;
  wire                _zz_435;
  wire       [1:0]    _zz_436;
  wire                _zz_437;
  wire       [1:0]    _zz_438;
  wire                _zz_439;
  wire       [1:0]    _zz_440;
  wire                _zz_441;
  wire       [1:0]    _zz_442;
  wire                _zz_443;
  wire       [1:0]    _zz_444;
  wire                _zz_445;
  wire       [1:0]    _zz_446;
  wire                _zz_447;
  wire       [1:0]    _zz_448;
  wire                _zz_449;
  wire       [1:0]    _zz_450;
  wire                _zz_451;
  wire       [1:0]    _zz_452;
  wire                _zz_453;
  wire       [1:0]    _zz_454;
  wire                _zz_455;
  wire       [1:0]    _zz_456;
  wire                _zz_457;
  wire       [1:0]    _zz_458;
  wire                _zz_459;
  wire                _zz_460;
  wire       [1:0]    _zz_461;
  wire                _zz_462;
  wire                _zz_463;
  wire       [1:0]    _zz_464;
  wire                _zz_465;
  wire                _zz_466;
  wire       [1:0]    _zz_467;
  wire                _zz_468;
  wire                _zz_469;
  wire       [1:0]    _zz_470;
  wire                _zz_471;
  wire                _zz_472;
  wire       [1:0]    _zz_473;
  wire                _zz_474;
  wire                _zz_475;
  wire       [1:0]    _zz_476;
  wire                _zz_477;
  wire                _zz_478;
  wire       [1:0]    _zz_479;
  wire                _zz_480;
  wire                _zz_481;
  wire       [1:0]    _zz_482;
  wire                _zz_483;
  wire                _zz_484;
  wire       [1:0]    _zz_485;
  wire                _zz_486;
  wire                _zz_487;
  wire       [1:0]    _zz_488;
  wire                _zz_489;
  wire                _zz_490;
  wire       [1:0]    _zz_491;
  wire                _zz_492;
  wire                _zz_493;
  wire       [1:0]    _zz_494;
  wire                _zz_495;
  wire                _zz_496;
  wire       [1:0]    _zz_497;
  wire                _zz_498;
  wire                _zz_499;
  wire       [1:0]    _zz_500;
  wire                _zz_501;
  wire                _zz_502;
  wire       [1:0]    _zz_503;
  wire                _zz_504;
  wire                _zz_505;
  wire       [1:0]    _zz_506;
  wire                _zz_507;
  wire                _zz_508;
  wire       [1:0]    _zz_509;
  wire                _zz_510;
  wire                _zz_511;
  wire       [1:0]    _zz_512;
  wire                _zz_513;
  wire                _zz_514;
  wire       [1:0]    _zz_515;
  wire                _zz_516;
  wire                _zz_517;
  wire       [1:0]    _zz_518;
  wire                _zz_519;
  wire                _zz_520;
  wire       [1:0]    _zz_521;
  wire                _zz_522;
  wire                _zz_523;
  wire       [1:0]    _zz_524;
  wire                _zz_525;
  wire                _zz_526;
  wire       [1:0]    _zz_527;
  wire                _zz_528;
  wire                _zz_529;
  wire       [1:0]    _zz_530;
  wire                _zz_531;
  wire                _zz_532;
  wire       [1:0]    _zz_533;
  wire                _zz_534;
  wire                _zz_535;
  wire       [1:0]    _zz_536;
  wire                _zz_537;
  wire                _zz_538;
  wire       [1:0]    _zz_539;
  wire                _zz_540;
  wire       [1:0]    _zz_541;
  wire                _zz_542;
  wire                _zz_543;
  wire       [1:0]    _zz_544;
  wire                _zz_545;
  wire                _zz_546;
  wire       [1:0]    _zz_547;
  wire                _zz_548;
  wire                _zz_549;
  wire       [1:0]    _zz_550;
  wire                _zz_551;
  wire                _zz_552;
  wire       [1:0]    _zz_553;
  wire                _zz_554;
  wire                _zz_555;
  wire       [1:0]    _zz_556;
  wire                _zz_557;
  wire                _zz_558;
  wire       [1:0]    _zz_559;
  wire                _zz_560;
  reg        [1:0]    _zz_561;
  reg        [6:0]    _zz_562;
  wire                _zz_563;
  wire       [6:0]    _zz_564;
  wire                bus_askWrite;
  wire                bus_askRead;
  wire                bus_doWrite;
  wire                bus_doRead;
  reg        [1:0]    _zz_565;
  reg        [1:0]    _zz_566;
  reg        [1:0]    _zz_567;
  reg        [1:0]    _zz_568;
  reg        [1:0]    _zz_569;
  reg        [1:0]    _zz_570;
  reg        [1:0]    _zz_571;
  reg        [1:0]    _zz_572;
  reg        [1:0]    _zz_573;
  reg        [1:0]    _zz_574;
  reg        [1:0]    _zz_575;
  reg        [1:0]    _zz_576;
  reg        [1:0]    _zz_577;
  reg        [1:0]    _zz_578;
  reg        [1:0]    _zz_579;
  reg        [1:0]    _zz_580;
  reg        [1:0]    _zz_581;
  reg        [1:0]    _zz_582;
  reg        [1:0]    _zz_583;
  reg        [1:0]    _zz_584;
  reg        [1:0]    _zz_585;
  reg        [1:0]    _zz_586;
  reg        [1:0]    _zz_587;
  reg        [1:0]    _zz_588;
  reg        [1:0]    _zz_589;
  reg        [1:0]    _zz_590;
  reg        [1:0]    _zz_591;
  reg        [1:0]    _zz_592;
  reg        [1:0]    _zz_593;
  reg        [1:0]    _zz_594;
  reg        [1:0]    _zz_595;
  reg        [1:0]    _zz_596;
  reg        [1:0]    _zz_597;
  reg        [1:0]    _zz_598;
  reg        [1:0]    _zz_599;
  reg                 mapping_claim_valid;
  reg        [6:0]    mapping_claim_payload;
  reg                 mapping_completion_valid;
  reg        [6:0]    mapping_completion_payload;
  reg                 mapping_coherencyStall_willIncrement;
  wire                mapping_coherencyStall_willClear;
  reg        [0:0]    mapping_coherencyStall_valueNext;
  reg        [0:0]    mapping_coherencyStall_value;
  wire                mapping_coherencyStall_willOverflowIfInc;
  wire                mapping_coherencyStall_willOverflow;
  reg        [1:0]    _zz_600;
  reg                 mapping_targetMapping_0_targetCompletion_valid;
  wire       [6:0]    mapping_targetMapping_0_targetCompletion_payload;
  reg                 _zz_601;
  reg                 _zz_602;
  reg                 _zz_603;
  reg                 _zz_604;
  reg                 _zz_605;
  reg                 _zz_606;
  reg                 _zz_607;
  reg                 _zz_608;
  reg                 _zz_609;
  reg                 _zz_610;
  reg                 _zz_611;
  reg                 _zz_612;
  reg                 _zz_613;
  reg                 _zz_614;
  reg                 _zz_615;
  reg                 _zz_616;
  reg                 _zz_617;
  reg                 _zz_618;
  reg                 _zz_619;
  reg                 _zz_620;
  reg                 _zz_621;
  reg                 _zz_622;
  reg                 _zz_623;
  reg                 _zz_624;
  reg                 _zz_625;
  reg                 _zz_626;
  reg                 _zz_627;
  reg                 _zz_628;
  reg                 _zz_629;
  reg                 _zz_630;
  reg                 _zz_631;
  reg                 _zz_632;
  reg                 _zz_633;
  reg                 _zz_634;
  reg                 _zz_635;
  reg        [1:0]    _zz_636;
  reg                 mapping_targetMapping_1_targetCompletion_valid;
  wire       [6:0]    mapping_targetMapping_1_targetCompletion_payload;
  reg                 _zz_637;
  reg                 _zz_638;
  reg                 _zz_639;
  reg                 _zz_640;
  reg                 _zz_641;
  reg                 _zz_642;
  reg                 _zz_643;
  reg                 _zz_644;
  reg                 _zz_645;
  reg                 _zz_646;
  reg                 _zz_647;
  reg                 _zz_648;
  reg                 _zz_649;
  reg                 _zz_650;
  reg                 _zz_651;
  reg                 _zz_652;
  reg                 _zz_653;
  reg                 _zz_654;
  reg                 _zz_655;
  reg                 _zz_656;
  reg                 _zz_657;
  reg                 _zz_658;
  reg                 _zz_659;
  reg                 _zz_660;
  reg                 _zz_661;
  reg                 _zz_662;
  reg                 _zz_663;
  reg                 _zz_664;
  reg                 _zz_665;
  reg                 _zz_666;
  reg                 _zz_667;
  reg                 _zz_668;
  reg                 _zz_669;
  reg                 _zz_670;
  reg                 _zz_671;
  reg        [1:0]    _zz_672;
  reg                 mapping_targetMapping_2_targetCompletion_valid;
  wire       [6:0]    mapping_targetMapping_2_targetCompletion_payload;
  reg                 _zz_673;
  reg                 _zz_674;
  reg                 _zz_675;
  reg                 _zz_676;
  reg                 _zz_677;
  reg                 _zz_678;
  reg                 _zz_679;
  reg                 _zz_680;
  reg                 _zz_681;
  reg                 _zz_682;
  reg                 _zz_683;
  reg                 _zz_684;
  reg                 _zz_685;
  reg                 _zz_686;
  reg                 _zz_687;
  reg                 _zz_688;
  reg                 _zz_689;
  reg                 _zz_690;
  reg                 _zz_691;
  reg                 _zz_692;
  reg                 _zz_693;
  reg                 _zz_694;
  reg                 _zz_695;
  reg                 _zz_696;
  reg                 _zz_697;
  reg                 _zz_698;
  reg                 _zz_699;
  reg                 _zz_700;
  reg                 _zz_701;
  reg                 _zz_702;
  reg                 _zz_703;
  reg                 _zz_704;
  reg                 _zz_705;
  reg                 _zz_706;
  reg                 _zz_707;

  assign _zz_708 = (mapping_coherencyStall_value != 1'b0);
  assign _zz_709 = io_apb_PWDATA[21 : 21];
  assign _zz_710 = io_apb_PWDATA[20 : 20];
  assign _zz_711 = io_apb_PWDATA[24 : 24];
  assign _zz_712 = io_apb_PWDATA[17 : 17];
  assign _zz_713 = io_apb_PWDATA[6 : 6];
  assign _zz_714 = io_apb_PWDATA[31 : 31];
  assign _zz_715 = io_apb_PWDATA[14 : 14];
  assign _zz_716 = io_apb_PWDATA[2 : 2];
  assign _zz_717 = io_apb_PWDATA[16 : 16];
  assign _zz_718 = io_apb_PWDATA[8 : 8];
  assign _zz_719 = io_apb_PWDATA[17 : 17];
  assign _zz_720 = io_apb_PWDATA[12 : 12];
  assign _zz_721 = io_apb_PWDATA[5 : 5];
  assign _zz_722 = io_apb_PWDATA[0 : 0];
  assign _zz_723 = io_apb_PWDATA[21 : 21];
  assign _zz_724 = io_apb_PWDATA[6 : 6];
  assign _zz_725 = io_apb_PWDATA[20 : 20];
  assign _zz_726 = io_apb_PWDATA[9 : 9];
  assign _zz_727 = io_apb_PWDATA[24 : 24];
  assign _zz_728 = io_apb_PWDATA[3 : 3];
  assign _zz_729 = io_apb_PWDATA[27 : 27];
  assign _zz_730 = io_apb_PWDATA[31 : 31];
  assign _zz_731 = io_apb_PWDATA[21 : 21];
  assign _zz_732 = io_apb_PWDATA[11 : 11];
  assign _zz_733 = io_apb_PWDATA[24 : 24];
  assign _zz_734 = io_apb_PWDATA[18 : 18];
  assign _zz_735 = io_apb_PWDATA[13 : 13];
  assign _zz_736 = io_apb_PWDATA[27 : 27];
  assign _zz_737 = io_apb_PWDATA[15 : 15];
  assign _zz_738 = io_apb_PWDATA[12 : 12];
  assign _zz_739 = io_apb_PWDATA[9 : 9];
  assign _zz_740 = io_apb_PWDATA[10 : 10];
  assign _zz_741 = io_apb_PWDATA[16 : 16];
  assign _zz_742 = io_apb_PWDATA[28 : 28];
  assign _zz_743 = io_apb_PWDATA[3 : 3];
  assign _zz_744 = io_apb_PWDATA[21 : 21];
  assign _zz_745 = io_apb_PWDATA[20 : 20];
  assign _zz_746 = io_apb_PWDATA[24 : 24];
  assign _zz_747 = io_apb_PWDATA[17 : 17];
  assign _zz_748 = io_apb_PWDATA[6 : 6];
  assign _zz_749 = io_apb_PWDATA[31 : 31];
  assign _zz_750 = io_apb_PWDATA[14 : 14];
  assign _zz_751 = io_apb_PWDATA[2 : 2];
  assign _zz_752 = io_apb_PWDATA[16 : 16];
  assign _zz_753 = io_apb_PWDATA[8 : 8];
  assign _zz_754 = io_apb_PWDATA[17 : 17];
  assign _zz_755 = io_apb_PWDATA[12 : 12];
  assign _zz_756 = io_apb_PWDATA[5 : 5];
  assign _zz_757 = io_apb_PWDATA[0 : 0];
  assign _zz_758 = io_apb_PWDATA[21 : 21];
  assign _zz_759 = io_apb_PWDATA[6 : 6];
  assign _zz_760 = io_apb_PWDATA[20 : 20];
  assign _zz_761 = io_apb_PWDATA[9 : 9];
  assign _zz_762 = io_apb_PWDATA[24 : 24];
  assign _zz_763 = io_apb_PWDATA[3 : 3];
  assign _zz_764 = io_apb_PWDATA[27 : 27];
  assign _zz_765 = io_apb_PWDATA[31 : 31];
  assign _zz_766 = io_apb_PWDATA[21 : 21];
  assign _zz_767 = io_apb_PWDATA[11 : 11];
  assign _zz_768 = io_apb_PWDATA[24 : 24];
  assign _zz_769 = io_apb_PWDATA[18 : 18];
  assign _zz_770 = io_apb_PWDATA[13 : 13];
  assign _zz_771 = io_apb_PWDATA[27 : 27];
  assign _zz_772 = io_apb_PWDATA[15 : 15];
  assign _zz_773 = io_apb_PWDATA[12 : 12];
  assign _zz_774 = io_apb_PWDATA[9 : 9];
  assign _zz_775 = io_apb_PWDATA[10 : 10];
  assign _zz_776 = io_apb_PWDATA[16 : 16];
  assign _zz_777 = io_apb_PWDATA[28 : 28];
  assign _zz_778 = io_apb_PWDATA[3 : 3];
  assign _zz_779 = io_apb_PWDATA[21 : 21];
  assign _zz_780 = io_apb_PWDATA[20 : 20];
  assign _zz_781 = io_apb_PWDATA[24 : 24];
  assign _zz_782 = io_apb_PWDATA[17 : 17];
  assign _zz_783 = io_apb_PWDATA[6 : 6];
  assign _zz_784 = io_apb_PWDATA[31 : 31];
  assign _zz_785 = io_apb_PWDATA[14 : 14];
  assign _zz_786 = io_apb_PWDATA[2 : 2];
  assign _zz_787 = io_apb_PWDATA[16 : 16];
  assign _zz_788 = io_apb_PWDATA[8 : 8];
  assign _zz_789 = io_apb_PWDATA[17 : 17];
  assign _zz_790 = io_apb_PWDATA[12 : 12];
  assign _zz_791 = io_apb_PWDATA[5 : 5];
  assign _zz_792 = io_apb_PWDATA[0 : 0];
  assign _zz_793 = io_apb_PWDATA[21 : 21];
  assign _zz_794 = io_apb_PWDATA[6 : 6];
  assign _zz_795 = io_apb_PWDATA[20 : 20];
  assign _zz_796 = io_apb_PWDATA[9 : 9];
  assign _zz_797 = io_apb_PWDATA[24 : 24];
  assign _zz_798 = io_apb_PWDATA[3 : 3];
  assign _zz_799 = io_apb_PWDATA[27 : 27];
  assign _zz_800 = io_apb_PWDATA[31 : 31];
  assign _zz_801 = io_apb_PWDATA[21 : 21];
  assign _zz_802 = io_apb_PWDATA[11 : 11];
  assign _zz_803 = io_apb_PWDATA[24 : 24];
  assign _zz_804 = io_apb_PWDATA[18 : 18];
  assign _zz_805 = io_apb_PWDATA[13 : 13];
  assign _zz_806 = io_apb_PWDATA[27 : 27];
  assign _zz_807 = io_apb_PWDATA[15 : 15];
  assign _zz_808 = io_apb_PWDATA[12 : 12];
  assign _zz_809 = io_apb_PWDATA[9 : 9];
  assign _zz_810 = io_apb_PWDATA[10 : 10];
  assign _zz_811 = io_apb_PWDATA[16 : 16];
  assign _zz_812 = io_apb_PWDATA[28 : 28];
  assign _zz_813 = io_apb_PWDATA[3 : 3];
  assign _zz_814 = (_zz_90 ? (_zz_36 ? targets_0_requests_0_id : targets_0_requests_1_id) : (_zz_39 ? targets_0_requests_2_id : targets_0_requests_3_id));
  assign _zz_815 = (_zz_93 ? (_zz_42 ? targets_0_requests_4_id : targets_0_requests_5_id) : (_zz_45 ? targets_0_requests_6_id : targets_0_requests_7_id));
  assign _zz_816 = (_zz_96 ? (_zz_48 ? targets_0_requests_8_id : targets_0_requests_9_id) : (_zz_51 ? targets_0_requests_10_id : targets_0_requests_11_id));
  assign _zz_817 = (_zz_99 ? (_zz_54 ? targets_0_requests_12_id : targets_0_requests_13_id) : (_zz_57 ? targets_0_requests_14_id : targets_0_requests_15_id));
  assign _zz_818 = (_zz_102 ? (_zz_60 ? targets_0_requests_16_id : targets_0_requests_17_id) : (_zz_63 ? targets_0_requests_18_id : targets_0_requests_19_id));
  assign _zz_819 = (_zz_105 ? (_zz_66 ? targets_0_requests_20_id : targets_0_requests_21_id) : (_zz_69 ? targets_0_requests_22_id : targets_0_requests_23_id));
  assign _zz_820 = (_zz_108 ? (_zz_72 ? targets_0_requests_24_id : targets_0_requests_25_id) : (_zz_75 ? targets_0_requests_26_id : targets_0_requests_27_id));
  assign _zz_821 = (_zz_111 ? (_zz_78 ? targets_0_requests_28_id : targets_0_requests_29_id) : (_zz_81 ? targets_0_requests_30_id : targets_0_requests_31_id));
  assign _zz_822 = (_zz_301 ? (_zz_247 ? _zz_830 : _zz_831) : (_zz_250 ? _zz_832 : _zz_833));
  assign _zz_823 = (_zz_304 ? (_zz_253 ? _zz_834 : _zz_835) : (_zz_256 ? _zz_836 : _zz_837));
  assign _zz_824 = (_zz_307 ? (_zz_259 ? _zz_838 : _zz_839) : (_zz_262 ? _zz_840 : _zz_841));
  assign _zz_825 = (_zz_310 ? (_zz_265 ? _zz_842 : _zz_843) : (_zz_268 ? _zz_844 : _zz_845));
  assign _zz_826 = (_zz_313 ? (_zz_271 ? _zz_846 : _zz_847) : (_zz_274 ? _zz_848 : _zz_849));
  assign _zz_827 = (_zz_316 ? (_zz_277 ? _zz_850 : _zz_851) : (_zz_280 ? _zz_852 : _zz_853));
  assign _zz_828 = (_zz_319 ? (_zz_283 ? _zz_854 : _zz_855) : (_zz_286 ? _zz_856 : _zz_857));
  assign _zz_829 = (_zz_322 ? (_zz_289 ? _zz_858 : _zz_859) : (_zz_292 ? _zz_860 : _zz_861));
  assign _zz_830 = 7'h0;
  assign _zz_831 = 7'h03;
  assign _zz_832 = 7'h0b;
  assign _zz_833 = 7'h12;
  assign _zz_834 = 7'h15;
  assign _zz_835 = 7'h18;
  assign _zz_836 = 7'h1b;
  assign _zz_837 = 7'h1f;
  assign _zz_838 = 7'h26;
  assign _zz_839 = 7'h31;
  assign _zz_840 = 7'h34;
  assign _zz_841 = 7'h35;
  assign _zz_842 = 7'h38;
  assign _zz_843 = 7'h3f;
  assign _zz_844 = 7'h40;
  assign _zz_845 = 7'h42;
  assign _zz_846 = 7'h45;
  assign _zz_847 = 7'h46;
  assign _zz_848 = 7'h48;
  assign _zz_849 = 7'h49;
  assign _zz_850 = 7'h4c;
  assign _zz_851 = 7'h4e;
  assign _zz_852 = 7'h50;
  assign _zz_853 = 7'h51;
  assign _zz_854 = 7'h54;
  assign _zz_855 = 7'h55;
  assign _zz_856 = 7'h58;
  assign _zz_857 = 7'h63;
  assign _zz_858 = 7'h69;
  assign _zz_859 = 7'h6a;
  assign _zz_860 = 7'h6c;
  assign _zz_861 = 7'h6d;
  assign _zz_862 = (_zz_514 ? (_zz_460 ? _zz_870 : _zz_871) : (_zz_463 ? _zz_872 : _zz_873));
  assign _zz_863 = (_zz_517 ? (_zz_466 ? _zz_874 : _zz_875) : (_zz_469 ? _zz_876 : _zz_877));
  assign _zz_864 = (_zz_520 ? (_zz_472 ? _zz_878 : _zz_879) : (_zz_475 ? _zz_880 : _zz_881));
  assign _zz_865 = (_zz_523 ? (_zz_478 ? _zz_882 : _zz_883) : (_zz_481 ? _zz_884 : _zz_885));
  assign _zz_866 = (_zz_526 ? (_zz_484 ? _zz_886 : _zz_887) : (_zz_487 ? _zz_888 : _zz_889));
  assign _zz_867 = (_zz_529 ? (_zz_490 ? _zz_890 : _zz_891) : (_zz_493 ? _zz_892 : _zz_893));
  assign _zz_868 = (_zz_532 ? (_zz_496 ? _zz_894 : _zz_895) : (_zz_499 ? _zz_896 : _zz_897));
  assign _zz_869 = (_zz_535 ? (_zz_502 ? _zz_898 : _zz_899) : (_zz_505 ? _zz_900 : _zz_901));
  assign _zz_870 = 7'h0;
  assign _zz_871 = 7'h03;
  assign _zz_872 = 7'h0b;
  assign _zz_873 = 7'h12;
  assign _zz_874 = 7'h15;
  assign _zz_875 = 7'h18;
  assign _zz_876 = 7'h1b;
  assign _zz_877 = 7'h1f;
  assign _zz_878 = 7'h26;
  assign _zz_879 = 7'h31;
  assign _zz_880 = 7'h34;
  assign _zz_881 = 7'h35;
  assign _zz_882 = 7'h38;
  assign _zz_883 = 7'h3f;
  assign _zz_884 = 7'h40;
  assign _zz_885 = 7'h42;
  assign _zz_886 = 7'h45;
  assign _zz_887 = 7'h46;
  assign _zz_888 = 7'h48;
  assign _zz_889 = 7'h49;
  assign _zz_890 = 7'h4c;
  assign _zz_891 = 7'h4e;
  assign _zz_892 = 7'h50;
  assign _zz_893 = 7'h51;
  assign _zz_894 = 7'h54;
  assign _zz_895 = 7'h55;
  assign _zz_896 = 7'h58;
  assign _zz_897 = 7'h63;
  assign _zz_898 = 7'h69;
  assign _zz_899 = 7'h6a;
  assign _zz_900 = 7'h6c;
  assign _zz_901 = 7'h6d;
  assign _zz_1 = io_sources[0];
  assign _zz_2 = io_sources[1];
  assign _zz_3 = io_sources[2];
  assign _zz_4 = io_sources[3];
  assign _zz_5 = io_sources[4];
  assign _zz_6 = io_sources[5];
  assign _zz_7 = io_sources[6];
  assign _zz_8 = io_sources[7];
  assign _zz_9 = io_sources[8];
  assign _zz_10 = io_sources[9];
  assign _zz_11 = io_sources[10];
  assign _zz_12 = io_sources[11];
  assign _zz_13 = io_sources[12];
  assign _zz_14 = io_sources[13];
  assign _zz_15 = io_sources[14];
  assign _zz_16 = io_sources[15];
  assign _zz_17 = io_sources[16];
  assign _zz_18 = io_sources[17];
  assign _zz_19 = io_sources[18];
  assign _zz_20 = io_sources[19];
  assign _zz_21 = io_sources[20];
  assign _zz_22 = io_sources[21];
  assign _zz_23 = io_sources[22];
  assign _zz_24 = io_sources[23];
  assign _zz_25 = io_sources[24];
  assign _zz_26 = io_sources[25];
  assign _zz_27 = io_sources[26];
  assign _zz_28 = io_sources[27];
  assign _zz_29 = io_sources[28];
  assign _zz_30 = io_sources[29];
  assign _zz_31 = io_sources[30];
  assign _zz_32 = io_sources[31];
  assign _zz_33 = io_sources[32];
  assign _zz_34 = io_sources[33];
  assign _zz_35 = io_sources[34];
  assign targets_0_requests_0_priority = 2'b00;
  assign targets_0_requests_0_id = 7'h0;
  assign targets_0_requests_0_valid = 1'b1;
  assign targets_0_requests_1_priority = gateways_2_priority;
  assign targets_0_requests_1_id = 7'h03;
  assign targets_0_requests_1_valid = (gateways_2_ip && targets_0_ie_2);
  assign targets_0_requests_2_priority = gateways_20_priority;
  assign targets_0_requests_2_id = 7'h0b;
  assign targets_0_requests_2_valid = (gateways_20_ip && targets_0_ie_20);
  assign targets_0_requests_3_priority = gateways_32_priority;
  assign targets_0_requests_3_id = 7'h12;
  assign targets_0_requests_3_valid = (gateways_32_ip && targets_0_ie_32);
  assign targets_0_requests_4_priority = gateways_15_priority;
  assign targets_0_requests_4_id = 7'h15;
  assign targets_0_requests_4_valid = (gateways_15_ip && targets_0_ie_15);
  assign targets_0_requests_5_priority = gateways_29_priority;
  assign targets_0_requests_5_id = 7'h18;
  assign targets_0_requests_5_valid = (gateways_29_ip && targets_0_ie_29);
  assign targets_0_requests_6_priority = gateways_3_priority;
  assign targets_0_requests_6_id = 7'h1b;
  assign targets_0_requests_6_valid = (gateways_3_ip && targets_0_ie_3);
  assign targets_0_requests_7_priority = gateways_7_priority;
  assign targets_0_requests_7_id = 7'h1f;
  assign targets_0_requests_7_valid = (gateways_7_ip && targets_0_ie_7);
  assign targets_0_requests_8_priority = gateways_24_priority;
  assign targets_0_requests_8_id = 7'h26;
  assign targets_0_requests_8_valid = (gateways_24_ip && targets_0_ie_24);
  assign targets_0_requests_9_priority = gateways_23_priority;
  assign targets_0_requests_9_id = 7'h31;
  assign targets_0_requests_9_valid = (gateways_23_ip && targets_0_ie_23);
  assign targets_0_requests_10_priority = gateways_14_priority;
  assign targets_0_requests_10_id = 7'h34;
  assign targets_0_requests_10_valid = (gateways_14_ip && targets_0_ie_14);
  assign targets_0_requests_11_priority = gateways_0_priority;
  assign targets_0_requests_11_id = 7'h35;
  assign targets_0_requests_11_valid = (gateways_0_ip && targets_0_ie_0);
  assign targets_0_requests_12_priority = gateways_21_priority;
  assign targets_0_requests_12_id = 7'h38;
  assign targets_0_requests_12_valid = (gateways_21_ip && targets_0_ie_21);
  assign targets_0_requests_13_priority = gateways_25_priority;
  assign targets_0_requests_13_id = 7'h3f;
  assign targets_0_requests_13_valid = (gateways_25_ip && targets_0_ie_25);
  assign targets_0_requests_14_priority = gateways_17_priority;
  assign targets_0_requests_14_id = 7'h40;
  assign targets_0_requests_14_valid = (gateways_17_ip && targets_0_ie_17);
  assign targets_0_requests_15_priority = gateways_5_priority;
  assign targets_0_requests_15_id = 7'h42;
  assign targets_0_requests_15_valid = (gateways_5_ip && targets_0_ie_5);
  assign targets_0_requests_16_priority = gateways_16_priority;
  assign targets_0_requests_16_id = 7'h45;
  assign targets_0_requests_16_valid = (gateways_16_ip && targets_0_ie_16);
  assign targets_0_requests_17_priority = gateways_22_priority;
  assign targets_0_requests_17_id = 7'h46;
  assign targets_0_requests_17_valid = (gateways_22_ip && targets_0_ie_22);
  assign targets_0_requests_18_priority = gateways_10_priority;
  assign targets_0_requests_18_id = 7'h48;
  assign targets_0_requests_18_valid = (gateways_10_ip && targets_0_ie_10);
  assign targets_0_requests_19_priority = gateways_31_priority;
  assign targets_0_requests_19_id = 7'h49;
  assign targets_0_requests_19_valid = (gateways_31_ip && targets_0_ie_31);
  assign targets_0_requests_20_priority = gateways_12_priority;
  assign targets_0_requests_20_id = 7'h4c;
  assign targets_0_requests_20_valid = (gateways_12_ip && targets_0_ie_12);
  assign targets_0_requests_21_priority = gateways_1_priority;
  assign targets_0_requests_21_id = 7'h4e;
  assign targets_0_requests_21_valid = (gateways_1_ip && targets_0_ie_1);
  assign targets_0_requests_22_priority = gateways_6_priority;
  assign targets_0_requests_22_id = 7'h50;
  assign targets_0_requests_22_valid = (gateways_6_ip && targets_0_ie_6);
  assign targets_0_requests_23_priority = gateways_11_priority;
  assign targets_0_requests_23_id = 7'h51;
  assign targets_0_requests_23_valid = (gateways_11_ip && targets_0_ie_11);
  assign targets_0_requests_24_priority = gateways_27_priority;
  assign targets_0_requests_24_id = 7'h54;
  assign targets_0_requests_24_valid = (gateways_27_ip && targets_0_ie_27);
  assign targets_0_requests_25_priority = gateways_19_priority;
  assign targets_0_requests_25_id = 7'h55;
  assign targets_0_requests_25_valid = (gateways_19_ip && targets_0_ie_19);
  assign targets_0_requests_26_priority = gateways_34_priority;
  assign targets_0_requests_26_id = 7'h58;
  assign targets_0_requests_26_valid = (gateways_34_ip && targets_0_ie_34);
  assign targets_0_requests_27_priority = gateways_33_priority;
  assign targets_0_requests_27_id = 7'h63;
  assign targets_0_requests_27_valid = (gateways_33_ip && targets_0_ie_33);
  assign targets_0_requests_28_priority = gateways_18_priority;
  assign targets_0_requests_28_id = 7'h69;
  assign targets_0_requests_28_valid = (gateways_18_ip && targets_0_ie_18);
  assign targets_0_requests_29_priority = gateways_26_priority;
  assign targets_0_requests_29_id = 7'h6a;
  assign targets_0_requests_29_valid = (gateways_26_ip && targets_0_ie_26);
  assign targets_0_requests_30_priority = gateways_13_priority;
  assign targets_0_requests_30_id = 7'h6c;
  assign targets_0_requests_30_valid = (gateways_13_ip && targets_0_ie_13);
  assign targets_0_requests_31_priority = gateways_4_priority;
  assign targets_0_requests_31_id = 7'h6d;
  assign targets_0_requests_31_valid = (gateways_4_ip && targets_0_ie_4);
  assign targets_0_requests_32_priority = gateways_9_priority;
  assign targets_0_requests_32_id = 7'h6f;
  assign targets_0_requests_32_valid = (gateways_9_ip && targets_0_ie_9);
  assign targets_0_requests_33_priority = gateways_28_priority;
  assign targets_0_requests_33_id = 7'h70;
  assign targets_0_requests_33_valid = (gateways_28_ip && targets_0_ie_28);
  assign targets_0_requests_34_priority = gateways_8_priority;
  assign targets_0_requests_34_id = 7'h7b;
  assign targets_0_requests_34_valid = (gateways_8_ip && targets_0_ie_8);
  assign targets_0_requests_35_priority = gateways_30_priority;
  assign targets_0_requests_35_id = 7'h7c;
  assign targets_0_requests_35_valid = (gateways_30_ip && targets_0_ie_30);
  assign _zz_36 = ((! targets_0_requests_1_valid) || (targets_0_requests_0_valid && (targets_0_requests_1_priority <= targets_0_requests_0_priority)));
  assign _zz_37 = (_zz_36 ? targets_0_requests_0_priority : targets_0_requests_1_priority);
  assign _zz_38 = (_zz_36 ? targets_0_requests_0_valid : targets_0_requests_1_valid);
  assign _zz_39 = ((! targets_0_requests_3_valid) || (targets_0_requests_2_valid && (targets_0_requests_3_priority <= targets_0_requests_2_priority)));
  assign _zz_40 = (_zz_39 ? targets_0_requests_2_priority : targets_0_requests_3_priority);
  assign _zz_41 = (_zz_39 ? targets_0_requests_2_valid : targets_0_requests_3_valid);
  assign _zz_42 = ((! targets_0_requests_5_valid) || (targets_0_requests_4_valid && (targets_0_requests_5_priority <= targets_0_requests_4_priority)));
  assign _zz_43 = (_zz_42 ? targets_0_requests_4_priority : targets_0_requests_5_priority);
  assign _zz_44 = (_zz_42 ? targets_0_requests_4_valid : targets_0_requests_5_valid);
  assign _zz_45 = ((! targets_0_requests_7_valid) || (targets_0_requests_6_valid && (targets_0_requests_7_priority <= targets_0_requests_6_priority)));
  assign _zz_46 = (_zz_45 ? targets_0_requests_6_priority : targets_0_requests_7_priority);
  assign _zz_47 = (_zz_45 ? targets_0_requests_6_valid : targets_0_requests_7_valid);
  assign _zz_48 = ((! targets_0_requests_9_valid) || (targets_0_requests_8_valid && (targets_0_requests_9_priority <= targets_0_requests_8_priority)));
  assign _zz_49 = (_zz_48 ? targets_0_requests_8_priority : targets_0_requests_9_priority);
  assign _zz_50 = (_zz_48 ? targets_0_requests_8_valid : targets_0_requests_9_valid);
  assign _zz_51 = ((! targets_0_requests_11_valid) || (targets_0_requests_10_valid && (targets_0_requests_11_priority <= targets_0_requests_10_priority)));
  assign _zz_52 = (_zz_51 ? targets_0_requests_10_priority : targets_0_requests_11_priority);
  assign _zz_53 = (_zz_51 ? targets_0_requests_10_valid : targets_0_requests_11_valid);
  assign _zz_54 = ((! targets_0_requests_13_valid) || (targets_0_requests_12_valid && (targets_0_requests_13_priority <= targets_0_requests_12_priority)));
  assign _zz_55 = (_zz_54 ? targets_0_requests_12_priority : targets_0_requests_13_priority);
  assign _zz_56 = (_zz_54 ? targets_0_requests_12_valid : targets_0_requests_13_valid);
  assign _zz_57 = ((! targets_0_requests_15_valid) || (targets_0_requests_14_valid && (targets_0_requests_15_priority <= targets_0_requests_14_priority)));
  assign _zz_58 = (_zz_57 ? targets_0_requests_14_priority : targets_0_requests_15_priority);
  assign _zz_59 = (_zz_57 ? targets_0_requests_14_valid : targets_0_requests_15_valid);
  assign _zz_60 = ((! targets_0_requests_17_valid) || (targets_0_requests_16_valid && (targets_0_requests_17_priority <= targets_0_requests_16_priority)));
  assign _zz_61 = (_zz_60 ? targets_0_requests_16_priority : targets_0_requests_17_priority);
  assign _zz_62 = (_zz_60 ? targets_0_requests_16_valid : targets_0_requests_17_valid);
  assign _zz_63 = ((! targets_0_requests_19_valid) || (targets_0_requests_18_valid && (targets_0_requests_19_priority <= targets_0_requests_18_priority)));
  assign _zz_64 = (_zz_63 ? targets_0_requests_18_priority : targets_0_requests_19_priority);
  assign _zz_65 = (_zz_63 ? targets_0_requests_18_valid : targets_0_requests_19_valid);
  assign _zz_66 = ((! targets_0_requests_21_valid) || (targets_0_requests_20_valid && (targets_0_requests_21_priority <= targets_0_requests_20_priority)));
  assign _zz_67 = (_zz_66 ? targets_0_requests_20_priority : targets_0_requests_21_priority);
  assign _zz_68 = (_zz_66 ? targets_0_requests_20_valid : targets_0_requests_21_valid);
  assign _zz_69 = ((! targets_0_requests_23_valid) || (targets_0_requests_22_valid && (targets_0_requests_23_priority <= targets_0_requests_22_priority)));
  assign _zz_70 = (_zz_69 ? targets_0_requests_22_priority : targets_0_requests_23_priority);
  assign _zz_71 = (_zz_69 ? targets_0_requests_22_valid : targets_0_requests_23_valid);
  assign _zz_72 = ((! targets_0_requests_25_valid) || (targets_0_requests_24_valid && (targets_0_requests_25_priority <= targets_0_requests_24_priority)));
  assign _zz_73 = (_zz_72 ? targets_0_requests_24_priority : targets_0_requests_25_priority);
  assign _zz_74 = (_zz_72 ? targets_0_requests_24_valid : targets_0_requests_25_valid);
  assign _zz_75 = ((! targets_0_requests_27_valid) || (targets_0_requests_26_valid && (targets_0_requests_27_priority <= targets_0_requests_26_priority)));
  assign _zz_76 = (_zz_75 ? targets_0_requests_26_priority : targets_0_requests_27_priority);
  assign _zz_77 = (_zz_75 ? targets_0_requests_26_valid : targets_0_requests_27_valid);
  assign _zz_78 = ((! targets_0_requests_29_valid) || (targets_0_requests_28_valid && (targets_0_requests_29_priority <= targets_0_requests_28_priority)));
  assign _zz_79 = (_zz_78 ? targets_0_requests_28_priority : targets_0_requests_29_priority);
  assign _zz_80 = (_zz_78 ? targets_0_requests_28_valid : targets_0_requests_29_valid);
  assign _zz_81 = ((! targets_0_requests_31_valid) || (targets_0_requests_30_valid && (targets_0_requests_31_priority <= targets_0_requests_30_priority)));
  assign _zz_82 = (_zz_81 ? targets_0_requests_30_priority : targets_0_requests_31_priority);
  assign _zz_83 = (_zz_81 ? targets_0_requests_30_valid : targets_0_requests_31_valid);
  assign _zz_84 = ((! targets_0_requests_33_valid) || (targets_0_requests_32_valid && (targets_0_requests_33_priority <= targets_0_requests_32_priority)));
  assign _zz_85 = (_zz_84 ? targets_0_requests_32_priority : targets_0_requests_33_priority);
  assign _zz_86 = (_zz_84 ? targets_0_requests_32_valid : targets_0_requests_33_valid);
  assign _zz_87 = ((! targets_0_requests_35_valid) || (targets_0_requests_34_valid && (targets_0_requests_35_priority <= targets_0_requests_34_priority)));
  assign _zz_88 = (_zz_87 ? targets_0_requests_34_priority : targets_0_requests_35_priority);
  assign _zz_89 = (_zz_87 ? targets_0_requests_34_valid : targets_0_requests_35_valid);
  assign _zz_90 = ((! _zz_41) || (_zz_38 && (_zz_40 <= _zz_37)));
  assign _zz_91 = (_zz_90 ? _zz_37 : _zz_40);
  assign _zz_92 = (_zz_90 ? _zz_38 : _zz_41);
  assign _zz_93 = ((! _zz_47) || (_zz_44 && (_zz_46 <= _zz_43)));
  assign _zz_94 = (_zz_93 ? _zz_43 : _zz_46);
  assign _zz_95 = (_zz_93 ? _zz_44 : _zz_47);
  assign _zz_96 = ((! _zz_53) || (_zz_50 && (_zz_52 <= _zz_49)));
  assign _zz_97 = (_zz_96 ? _zz_49 : _zz_52);
  assign _zz_98 = (_zz_96 ? _zz_50 : _zz_53);
  assign _zz_99 = ((! _zz_59) || (_zz_56 && (_zz_58 <= _zz_55)));
  assign _zz_100 = (_zz_99 ? _zz_55 : _zz_58);
  assign _zz_101 = (_zz_99 ? _zz_56 : _zz_59);
  assign _zz_102 = ((! _zz_65) || (_zz_62 && (_zz_64 <= _zz_61)));
  assign _zz_103 = (_zz_102 ? _zz_61 : _zz_64);
  assign _zz_104 = (_zz_102 ? _zz_62 : _zz_65);
  assign _zz_105 = ((! _zz_71) || (_zz_68 && (_zz_70 <= _zz_67)));
  assign _zz_106 = (_zz_105 ? _zz_67 : _zz_70);
  assign _zz_107 = (_zz_105 ? _zz_68 : _zz_71);
  assign _zz_108 = ((! _zz_77) || (_zz_74 && (_zz_76 <= _zz_73)));
  assign _zz_109 = (_zz_108 ? _zz_73 : _zz_76);
  assign _zz_110 = (_zz_108 ? _zz_74 : _zz_77);
  assign _zz_111 = ((! _zz_83) || (_zz_80 && (_zz_82 <= _zz_79)));
  assign _zz_112 = (_zz_111 ? _zz_79 : _zz_82);
  assign _zz_113 = (_zz_111 ? _zz_80 : _zz_83);
  assign _zz_114 = ((! _zz_89) || (_zz_86 && (_zz_88 <= _zz_85)));
  assign _zz_115 = (_zz_114 ? _zz_85 : _zz_88);
  assign _zz_116 = (_zz_114 ? _zz_86 : _zz_89);
  assign _zz_117 = ((! _zz_95) || (_zz_92 && (_zz_94 <= _zz_91)));
  assign _zz_118 = (_zz_117 ? _zz_91 : _zz_94);
  assign _zz_119 = (_zz_117 ? _zz_92 : _zz_95);
  assign _zz_120 = ((! _zz_101) || (_zz_98 && (_zz_100 <= _zz_97)));
  assign _zz_121 = (_zz_120 ? _zz_97 : _zz_100);
  assign _zz_122 = (_zz_120 ? _zz_98 : _zz_101);
  assign _zz_123 = ((! _zz_107) || (_zz_104 && (_zz_106 <= _zz_103)));
  assign _zz_124 = (_zz_123 ? _zz_103 : _zz_106);
  assign _zz_125 = (_zz_123 ? _zz_104 : _zz_107);
  assign _zz_126 = ((! _zz_113) || (_zz_110 && (_zz_112 <= _zz_109)));
  assign _zz_127 = (_zz_126 ? _zz_109 : _zz_112);
  assign _zz_128 = (_zz_126 ? _zz_110 : _zz_113);
  assign _zz_129 = ((! _zz_122) || (_zz_119 && (_zz_121 <= _zz_118)));
  assign _zz_130 = (_zz_129 ? _zz_118 : _zz_121);
  assign _zz_131 = (_zz_129 ? _zz_119 : _zz_122);
  assign _zz_132 = ((! _zz_128) || (_zz_125 && (_zz_127 <= _zz_124)));
  assign _zz_133 = (_zz_132 ? _zz_124 : _zz_127);
  assign _zz_134 = (_zz_132 ? _zz_125 : _zz_128);
  assign _zz_135 = ((! _zz_134) || (_zz_131 && (_zz_133 <= _zz_130)));
  assign _zz_136 = (_zz_135 ? _zz_130 : _zz_133);
  assign _zz_137 = (_zz_135 ? _zz_131 : _zz_134);
  assign _zz_138 = ((! _zz_116) || (_zz_137 && (_zz_115 <= _zz_136)));
  assign targets_0_iep = (targets_0_threshold < targets_0_bestRequest_priority);
  assign targets_0_claim = (targets_0_iep ? targets_0_bestRequest_id : 7'h0);
  assign _zz_175 = 2'b00;
  assign _zz_176 = 1'b1;
  assign _zz_177 = gateways_2_priority;
  assign _zz_178 = (gateways_2_ip && _zz_141);
  assign _zz_179 = gateways_20_priority;
  assign _zz_180 = (gateways_20_ip && _zz_159);
  assign _zz_181 = gateways_32_priority;
  assign _zz_182 = (gateways_32_ip && _zz_171);
  assign _zz_183 = gateways_15_priority;
  assign _zz_184 = (gateways_15_ip && _zz_154);
  assign _zz_185 = gateways_29_priority;
  assign _zz_186 = (gateways_29_ip && _zz_168);
  assign _zz_187 = gateways_3_priority;
  assign _zz_188 = (gateways_3_ip && _zz_142);
  assign _zz_189 = gateways_7_priority;
  assign _zz_190 = (gateways_7_ip && _zz_146);
  assign _zz_191 = gateways_24_priority;
  assign _zz_192 = (gateways_24_ip && _zz_163);
  assign _zz_193 = gateways_23_priority;
  assign _zz_194 = (gateways_23_ip && _zz_162);
  assign _zz_195 = gateways_14_priority;
  assign _zz_196 = (gateways_14_ip && _zz_153);
  assign _zz_197 = gateways_0_priority;
  assign _zz_198 = (gateways_0_ip && _zz_139);
  assign _zz_199 = gateways_21_priority;
  assign _zz_200 = (gateways_21_ip && _zz_160);
  assign _zz_201 = gateways_25_priority;
  assign _zz_202 = (gateways_25_ip && _zz_164);
  assign _zz_203 = gateways_17_priority;
  assign _zz_204 = (gateways_17_ip && _zz_156);
  assign _zz_205 = gateways_5_priority;
  assign _zz_206 = (gateways_5_ip && _zz_144);
  assign _zz_207 = gateways_16_priority;
  assign _zz_208 = (gateways_16_ip && _zz_155);
  assign _zz_209 = gateways_22_priority;
  assign _zz_210 = (gateways_22_ip && _zz_161);
  assign _zz_211 = gateways_10_priority;
  assign _zz_212 = (gateways_10_ip && _zz_149);
  assign _zz_213 = gateways_31_priority;
  assign _zz_214 = (gateways_31_ip && _zz_170);
  assign _zz_215 = gateways_12_priority;
  assign _zz_216 = (gateways_12_ip && _zz_151);
  assign _zz_217 = gateways_1_priority;
  assign _zz_218 = (gateways_1_ip && _zz_140);
  assign _zz_219 = gateways_6_priority;
  assign _zz_220 = (gateways_6_ip && _zz_145);
  assign _zz_221 = gateways_11_priority;
  assign _zz_222 = (gateways_11_ip && _zz_150);
  assign _zz_223 = gateways_27_priority;
  assign _zz_224 = (gateways_27_ip && _zz_166);
  assign _zz_225 = gateways_19_priority;
  assign _zz_226 = (gateways_19_ip && _zz_158);
  assign _zz_227 = gateways_34_priority;
  assign _zz_228 = (gateways_34_ip && _zz_173);
  assign _zz_229 = gateways_33_priority;
  assign _zz_230 = (gateways_33_ip && _zz_172);
  assign _zz_231 = gateways_18_priority;
  assign _zz_232 = (gateways_18_ip && _zz_157);
  assign _zz_233 = gateways_26_priority;
  assign _zz_234 = (gateways_26_ip && _zz_165);
  assign _zz_235 = gateways_13_priority;
  assign _zz_236 = (gateways_13_ip && _zz_152);
  assign _zz_237 = gateways_4_priority;
  assign _zz_238 = (gateways_4_ip && _zz_143);
  assign _zz_239 = gateways_9_priority;
  assign _zz_240 = (gateways_9_ip && _zz_148);
  assign _zz_241 = gateways_28_priority;
  assign _zz_242 = (gateways_28_ip && _zz_167);
  assign _zz_243 = gateways_8_priority;
  assign _zz_244 = (gateways_8_ip && _zz_147);
  assign _zz_245 = gateways_30_priority;
  assign _zz_246 = (gateways_30_ip && _zz_169);
  assign _zz_247 = ((! _zz_178) || (_zz_176 && (_zz_177 <= _zz_175)));
  assign _zz_248 = (_zz_247 ? _zz_175 : _zz_177);
  assign _zz_249 = (_zz_247 ? _zz_176 : _zz_178);
  assign _zz_250 = ((! _zz_182) || (_zz_180 && (_zz_181 <= _zz_179)));
  assign _zz_251 = (_zz_250 ? _zz_179 : _zz_181);
  assign _zz_252 = (_zz_250 ? _zz_180 : _zz_182);
  assign _zz_253 = ((! _zz_186) || (_zz_184 && (_zz_185 <= _zz_183)));
  assign _zz_254 = (_zz_253 ? _zz_183 : _zz_185);
  assign _zz_255 = (_zz_253 ? _zz_184 : _zz_186);
  assign _zz_256 = ((! _zz_190) || (_zz_188 && (_zz_189 <= _zz_187)));
  assign _zz_257 = (_zz_256 ? _zz_187 : _zz_189);
  assign _zz_258 = (_zz_256 ? _zz_188 : _zz_190);
  assign _zz_259 = ((! _zz_194) || (_zz_192 && (_zz_193 <= _zz_191)));
  assign _zz_260 = (_zz_259 ? _zz_191 : _zz_193);
  assign _zz_261 = (_zz_259 ? _zz_192 : _zz_194);
  assign _zz_262 = ((! _zz_198) || (_zz_196 && (_zz_197 <= _zz_195)));
  assign _zz_263 = (_zz_262 ? _zz_195 : _zz_197);
  assign _zz_264 = (_zz_262 ? _zz_196 : _zz_198);
  assign _zz_265 = ((! _zz_202) || (_zz_200 && (_zz_201 <= _zz_199)));
  assign _zz_266 = (_zz_265 ? _zz_199 : _zz_201);
  assign _zz_267 = (_zz_265 ? _zz_200 : _zz_202);
  assign _zz_268 = ((! _zz_206) || (_zz_204 && (_zz_205 <= _zz_203)));
  assign _zz_269 = (_zz_268 ? _zz_203 : _zz_205);
  assign _zz_270 = (_zz_268 ? _zz_204 : _zz_206);
  assign _zz_271 = ((! _zz_210) || (_zz_208 && (_zz_209 <= _zz_207)));
  assign _zz_272 = (_zz_271 ? _zz_207 : _zz_209);
  assign _zz_273 = (_zz_271 ? _zz_208 : _zz_210);
  assign _zz_274 = ((! _zz_214) || (_zz_212 && (_zz_213 <= _zz_211)));
  assign _zz_275 = (_zz_274 ? _zz_211 : _zz_213);
  assign _zz_276 = (_zz_274 ? _zz_212 : _zz_214);
  assign _zz_277 = ((! _zz_218) || (_zz_216 && (_zz_217 <= _zz_215)));
  assign _zz_278 = (_zz_277 ? _zz_215 : _zz_217);
  assign _zz_279 = (_zz_277 ? _zz_216 : _zz_218);
  assign _zz_280 = ((! _zz_222) || (_zz_220 && (_zz_221 <= _zz_219)));
  assign _zz_281 = (_zz_280 ? _zz_219 : _zz_221);
  assign _zz_282 = (_zz_280 ? _zz_220 : _zz_222);
  assign _zz_283 = ((! _zz_226) || (_zz_224 && (_zz_225 <= _zz_223)));
  assign _zz_284 = (_zz_283 ? _zz_223 : _zz_225);
  assign _zz_285 = (_zz_283 ? _zz_224 : _zz_226);
  assign _zz_286 = ((! _zz_230) || (_zz_228 && (_zz_229 <= _zz_227)));
  assign _zz_287 = (_zz_286 ? _zz_227 : _zz_229);
  assign _zz_288 = (_zz_286 ? _zz_228 : _zz_230);
  assign _zz_289 = ((! _zz_234) || (_zz_232 && (_zz_233 <= _zz_231)));
  assign _zz_290 = (_zz_289 ? _zz_231 : _zz_233);
  assign _zz_291 = (_zz_289 ? _zz_232 : _zz_234);
  assign _zz_292 = ((! _zz_238) || (_zz_236 && (_zz_237 <= _zz_235)));
  assign _zz_293 = (_zz_292 ? _zz_235 : _zz_237);
  assign _zz_294 = (_zz_292 ? _zz_236 : _zz_238);
  assign _zz_295 = ((! _zz_242) || (_zz_240 && (_zz_241 <= _zz_239)));
  assign _zz_296 = (_zz_295 ? _zz_239 : _zz_241);
  assign _zz_297 = (_zz_295 ? _zz_240 : _zz_242);
  assign _zz_298 = ((! _zz_246) || (_zz_244 && (_zz_245 <= _zz_243)));
  assign _zz_299 = (_zz_298 ? _zz_243 : _zz_245);
  assign _zz_300 = (_zz_298 ? _zz_244 : _zz_246);
  assign _zz_301 = ((! _zz_252) || (_zz_249 && (_zz_251 <= _zz_248)));
  assign _zz_302 = (_zz_301 ? _zz_248 : _zz_251);
  assign _zz_303 = (_zz_301 ? _zz_249 : _zz_252);
  assign _zz_304 = ((! _zz_258) || (_zz_255 && (_zz_257 <= _zz_254)));
  assign _zz_305 = (_zz_304 ? _zz_254 : _zz_257);
  assign _zz_306 = (_zz_304 ? _zz_255 : _zz_258);
  assign _zz_307 = ((! _zz_264) || (_zz_261 && (_zz_263 <= _zz_260)));
  assign _zz_308 = (_zz_307 ? _zz_260 : _zz_263);
  assign _zz_309 = (_zz_307 ? _zz_261 : _zz_264);
  assign _zz_310 = ((! _zz_270) || (_zz_267 && (_zz_269 <= _zz_266)));
  assign _zz_311 = (_zz_310 ? _zz_266 : _zz_269);
  assign _zz_312 = (_zz_310 ? _zz_267 : _zz_270);
  assign _zz_313 = ((! _zz_276) || (_zz_273 && (_zz_275 <= _zz_272)));
  assign _zz_314 = (_zz_313 ? _zz_272 : _zz_275);
  assign _zz_315 = (_zz_313 ? _zz_273 : _zz_276);
  assign _zz_316 = ((! _zz_282) || (_zz_279 && (_zz_281 <= _zz_278)));
  assign _zz_317 = (_zz_316 ? _zz_278 : _zz_281);
  assign _zz_318 = (_zz_316 ? _zz_279 : _zz_282);
  assign _zz_319 = ((! _zz_288) || (_zz_285 && (_zz_287 <= _zz_284)));
  assign _zz_320 = (_zz_319 ? _zz_284 : _zz_287);
  assign _zz_321 = (_zz_319 ? _zz_285 : _zz_288);
  assign _zz_322 = ((! _zz_294) || (_zz_291 && (_zz_293 <= _zz_290)));
  assign _zz_323 = (_zz_322 ? _zz_290 : _zz_293);
  assign _zz_324 = (_zz_322 ? _zz_291 : _zz_294);
  assign _zz_325 = ((! _zz_300) || (_zz_297 && (_zz_299 <= _zz_296)));
  assign _zz_326 = (_zz_325 ? _zz_296 : _zz_299);
  assign _zz_327 = ((! _zz_306) || (_zz_303 && (_zz_305 <= _zz_302)));
  assign _zz_328 = (_zz_327 ? _zz_302 : _zz_305);
  assign _zz_329 = (_zz_327 ? _zz_303 : _zz_306);
  assign _zz_330 = ((! _zz_312) || (_zz_309 && (_zz_311 <= _zz_308)));
  assign _zz_331 = (_zz_330 ? _zz_308 : _zz_311);
  assign _zz_332 = (_zz_330 ? _zz_309 : _zz_312);
  assign _zz_333 = ((! _zz_318) || (_zz_315 && (_zz_317 <= _zz_314)));
  assign _zz_334 = (_zz_333 ? _zz_314 : _zz_317);
  assign _zz_335 = (_zz_333 ? _zz_315 : _zz_318);
  assign _zz_336 = ((! _zz_324) || (_zz_321 && (_zz_323 <= _zz_320)));
  assign _zz_337 = (_zz_336 ? _zz_320 : _zz_323);
  assign _zz_338 = (_zz_336 ? _zz_321 : _zz_324);
  assign _zz_339 = ((! _zz_332) || (_zz_329 && (_zz_331 <= _zz_328)));
  assign _zz_340 = (_zz_339 ? _zz_328 : _zz_331);
  assign _zz_341 = (_zz_339 ? _zz_329 : _zz_332);
  assign _zz_342 = ((! _zz_338) || (_zz_335 && (_zz_337 <= _zz_334)));
  assign _zz_343 = (_zz_342 ? _zz_334 : _zz_337);
  assign _zz_344 = (_zz_342 ? _zz_335 : _zz_338);
  assign _zz_345 = ((! _zz_344) || (_zz_341 && (_zz_343 <= _zz_340)));
  assign _zz_346 = (_zz_345 ? _zz_340 : _zz_343);
  assign _zz_347 = ((! (_zz_325 ? _zz_297 : _zz_300)) || ((_zz_345 ? _zz_341 : _zz_344) && (_zz_326 <= _zz_346)));
  assign _zz_350 = (_zz_174 < _zz_348);
  assign _zz_351 = (_zz_350 ? _zz_349 : 7'h0);
  assign _zz_388 = 2'b00;
  assign _zz_389 = 1'b1;
  assign _zz_390 = gateways_2_priority;
  assign _zz_391 = (gateways_2_ip && _zz_354);
  assign _zz_392 = gateways_20_priority;
  assign _zz_393 = (gateways_20_ip && _zz_372);
  assign _zz_394 = gateways_32_priority;
  assign _zz_395 = (gateways_32_ip && _zz_384);
  assign _zz_396 = gateways_15_priority;
  assign _zz_397 = (gateways_15_ip && _zz_367);
  assign _zz_398 = gateways_29_priority;
  assign _zz_399 = (gateways_29_ip && _zz_381);
  assign _zz_400 = gateways_3_priority;
  assign _zz_401 = (gateways_3_ip && _zz_355);
  assign _zz_402 = gateways_7_priority;
  assign _zz_403 = (gateways_7_ip && _zz_359);
  assign _zz_404 = gateways_24_priority;
  assign _zz_405 = (gateways_24_ip && _zz_376);
  assign _zz_406 = gateways_23_priority;
  assign _zz_407 = (gateways_23_ip && _zz_375);
  assign _zz_408 = gateways_14_priority;
  assign _zz_409 = (gateways_14_ip && _zz_366);
  assign _zz_410 = gateways_0_priority;
  assign _zz_411 = (gateways_0_ip && _zz_352);
  assign _zz_412 = gateways_21_priority;
  assign _zz_413 = (gateways_21_ip && _zz_373);
  assign _zz_414 = gateways_25_priority;
  assign _zz_415 = (gateways_25_ip && _zz_377);
  assign _zz_416 = gateways_17_priority;
  assign _zz_417 = (gateways_17_ip && _zz_369);
  assign _zz_418 = gateways_5_priority;
  assign _zz_419 = (gateways_5_ip && _zz_357);
  assign _zz_420 = gateways_16_priority;
  assign _zz_421 = (gateways_16_ip && _zz_368);
  assign _zz_422 = gateways_22_priority;
  assign _zz_423 = (gateways_22_ip && _zz_374);
  assign _zz_424 = gateways_10_priority;
  assign _zz_425 = (gateways_10_ip && _zz_362);
  assign _zz_426 = gateways_31_priority;
  assign _zz_427 = (gateways_31_ip && _zz_383);
  assign _zz_428 = gateways_12_priority;
  assign _zz_429 = (gateways_12_ip && _zz_364);
  assign _zz_430 = gateways_1_priority;
  assign _zz_431 = (gateways_1_ip && _zz_353);
  assign _zz_432 = gateways_6_priority;
  assign _zz_433 = (gateways_6_ip && _zz_358);
  assign _zz_434 = gateways_11_priority;
  assign _zz_435 = (gateways_11_ip && _zz_363);
  assign _zz_436 = gateways_27_priority;
  assign _zz_437 = (gateways_27_ip && _zz_379);
  assign _zz_438 = gateways_19_priority;
  assign _zz_439 = (gateways_19_ip && _zz_371);
  assign _zz_440 = gateways_34_priority;
  assign _zz_441 = (gateways_34_ip && _zz_386);
  assign _zz_442 = gateways_33_priority;
  assign _zz_443 = (gateways_33_ip && _zz_385);
  assign _zz_444 = gateways_18_priority;
  assign _zz_445 = (gateways_18_ip && _zz_370);
  assign _zz_446 = gateways_26_priority;
  assign _zz_447 = (gateways_26_ip && _zz_378);
  assign _zz_448 = gateways_13_priority;
  assign _zz_449 = (gateways_13_ip && _zz_365);
  assign _zz_450 = gateways_4_priority;
  assign _zz_451 = (gateways_4_ip && _zz_356);
  assign _zz_452 = gateways_9_priority;
  assign _zz_453 = (gateways_9_ip && _zz_361);
  assign _zz_454 = gateways_28_priority;
  assign _zz_455 = (gateways_28_ip && _zz_380);
  assign _zz_456 = gateways_8_priority;
  assign _zz_457 = (gateways_8_ip && _zz_360);
  assign _zz_458 = gateways_30_priority;
  assign _zz_459 = (gateways_30_ip && _zz_382);
  assign _zz_460 = ((! _zz_391) || (_zz_389 && (_zz_390 <= _zz_388)));
  assign _zz_461 = (_zz_460 ? _zz_388 : _zz_390);
  assign _zz_462 = (_zz_460 ? _zz_389 : _zz_391);
  assign _zz_463 = ((! _zz_395) || (_zz_393 && (_zz_394 <= _zz_392)));
  assign _zz_464 = (_zz_463 ? _zz_392 : _zz_394);
  assign _zz_465 = (_zz_463 ? _zz_393 : _zz_395);
  assign _zz_466 = ((! _zz_399) || (_zz_397 && (_zz_398 <= _zz_396)));
  assign _zz_467 = (_zz_466 ? _zz_396 : _zz_398);
  assign _zz_468 = (_zz_466 ? _zz_397 : _zz_399);
  assign _zz_469 = ((! _zz_403) || (_zz_401 && (_zz_402 <= _zz_400)));
  assign _zz_470 = (_zz_469 ? _zz_400 : _zz_402);
  assign _zz_471 = (_zz_469 ? _zz_401 : _zz_403);
  assign _zz_472 = ((! _zz_407) || (_zz_405 && (_zz_406 <= _zz_404)));
  assign _zz_473 = (_zz_472 ? _zz_404 : _zz_406);
  assign _zz_474 = (_zz_472 ? _zz_405 : _zz_407);
  assign _zz_475 = ((! _zz_411) || (_zz_409 && (_zz_410 <= _zz_408)));
  assign _zz_476 = (_zz_475 ? _zz_408 : _zz_410);
  assign _zz_477 = (_zz_475 ? _zz_409 : _zz_411);
  assign _zz_478 = ((! _zz_415) || (_zz_413 && (_zz_414 <= _zz_412)));
  assign _zz_479 = (_zz_478 ? _zz_412 : _zz_414);
  assign _zz_480 = (_zz_478 ? _zz_413 : _zz_415);
  assign _zz_481 = ((! _zz_419) || (_zz_417 && (_zz_418 <= _zz_416)));
  assign _zz_482 = (_zz_481 ? _zz_416 : _zz_418);
  assign _zz_483 = (_zz_481 ? _zz_417 : _zz_419);
  assign _zz_484 = ((! _zz_423) || (_zz_421 && (_zz_422 <= _zz_420)));
  assign _zz_485 = (_zz_484 ? _zz_420 : _zz_422);
  assign _zz_486 = (_zz_484 ? _zz_421 : _zz_423);
  assign _zz_487 = ((! _zz_427) || (_zz_425 && (_zz_426 <= _zz_424)));
  assign _zz_488 = (_zz_487 ? _zz_424 : _zz_426);
  assign _zz_489 = (_zz_487 ? _zz_425 : _zz_427);
  assign _zz_490 = ((! _zz_431) || (_zz_429 && (_zz_430 <= _zz_428)));
  assign _zz_491 = (_zz_490 ? _zz_428 : _zz_430);
  assign _zz_492 = (_zz_490 ? _zz_429 : _zz_431);
  assign _zz_493 = ((! _zz_435) || (_zz_433 && (_zz_434 <= _zz_432)));
  assign _zz_494 = (_zz_493 ? _zz_432 : _zz_434);
  assign _zz_495 = (_zz_493 ? _zz_433 : _zz_435);
  assign _zz_496 = ((! _zz_439) || (_zz_437 && (_zz_438 <= _zz_436)));
  assign _zz_497 = (_zz_496 ? _zz_436 : _zz_438);
  assign _zz_498 = (_zz_496 ? _zz_437 : _zz_439);
  assign _zz_499 = ((! _zz_443) || (_zz_441 && (_zz_442 <= _zz_440)));
  assign _zz_500 = (_zz_499 ? _zz_440 : _zz_442);
  assign _zz_501 = (_zz_499 ? _zz_441 : _zz_443);
  assign _zz_502 = ((! _zz_447) || (_zz_445 && (_zz_446 <= _zz_444)));
  assign _zz_503 = (_zz_502 ? _zz_444 : _zz_446);
  assign _zz_504 = (_zz_502 ? _zz_445 : _zz_447);
  assign _zz_505 = ((! _zz_451) || (_zz_449 && (_zz_450 <= _zz_448)));
  assign _zz_506 = (_zz_505 ? _zz_448 : _zz_450);
  assign _zz_507 = (_zz_505 ? _zz_449 : _zz_451);
  assign _zz_508 = ((! _zz_455) || (_zz_453 && (_zz_454 <= _zz_452)));
  assign _zz_509 = (_zz_508 ? _zz_452 : _zz_454);
  assign _zz_510 = (_zz_508 ? _zz_453 : _zz_455);
  assign _zz_511 = ((! _zz_459) || (_zz_457 && (_zz_458 <= _zz_456)));
  assign _zz_512 = (_zz_511 ? _zz_456 : _zz_458);
  assign _zz_513 = (_zz_511 ? _zz_457 : _zz_459);
  assign _zz_514 = ((! _zz_465) || (_zz_462 && (_zz_464 <= _zz_461)));
  assign _zz_515 = (_zz_514 ? _zz_461 : _zz_464);
  assign _zz_516 = (_zz_514 ? _zz_462 : _zz_465);
  assign _zz_517 = ((! _zz_471) || (_zz_468 && (_zz_470 <= _zz_467)));
  assign _zz_518 = (_zz_517 ? _zz_467 : _zz_470);
  assign _zz_519 = (_zz_517 ? _zz_468 : _zz_471);
  assign _zz_520 = ((! _zz_477) || (_zz_474 && (_zz_476 <= _zz_473)));
  assign _zz_521 = (_zz_520 ? _zz_473 : _zz_476);
  assign _zz_522 = (_zz_520 ? _zz_474 : _zz_477);
  assign _zz_523 = ((! _zz_483) || (_zz_480 && (_zz_482 <= _zz_479)));
  assign _zz_524 = (_zz_523 ? _zz_479 : _zz_482);
  assign _zz_525 = (_zz_523 ? _zz_480 : _zz_483);
  assign _zz_526 = ((! _zz_489) || (_zz_486 && (_zz_488 <= _zz_485)));
  assign _zz_527 = (_zz_526 ? _zz_485 : _zz_488);
  assign _zz_528 = (_zz_526 ? _zz_486 : _zz_489);
  assign _zz_529 = ((! _zz_495) || (_zz_492 && (_zz_494 <= _zz_491)));
  assign _zz_530 = (_zz_529 ? _zz_491 : _zz_494);
  assign _zz_531 = (_zz_529 ? _zz_492 : _zz_495);
  assign _zz_532 = ((! _zz_501) || (_zz_498 && (_zz_500 <= _zz_497)));
  assign _zz_533 = (_zz_532 ? _zz_497 : _zz_500);
  assign _zz_534 = (_zz_532 ? _zz_498 : _zz_501);
  assign _zz_535 = ((! _zz_507) || (_zz_504 && (_zz_506 <= _zz_503)));
  assign _zz_536 = (_zz_535 ? _zz_503 : _zz_506);
  assign _zz_537 = (_zz_535 ? _zz_504 : _zz_507);
  assign _zz_538 = ((! _zz_513) || (_zz_510 && (_zz_512 <= _zz_509)));
  assign _zz_539 = (_zz_538 ? _zz_509 : _zz_512);
  assign _zz_540 = ((! _zz_519) || (_zz_516 && (_zz_518 <= _zz_515)));
  assign _zz_541 = (_zz_540 ? _zz_515 : _zz_518);
  assign _zz_542 = (_zz_540 ? _zz_516 : _zz_519);
  assign _zz_543 = ((! _zz_525) || (_zz_522 && (_zz_524 <= _zz_521)));
  assign _zz_544 = (_zz_543 ? _zz_521 : _zz_524);
  assign _zz_545 = (_zz_543 ? _zz_522 : _zz_525);
  assign _zz_546 = ((! _zz_531) || (_zz_528 && (_zz_530 <= _zz_527)));
  assign _zz_547 = (_zz_546 ? _zz_527 : _zz_530);
  assign _zz_548 = (_zz_546 ? _zz_528 : _zz_531);
  assign _zz_549 = ((! _zz_537) || (_zz_534 && (_zz_536 <= _zz_533)));
  assign _zz_550 = (_zz_549 ? _zz_533 : _zz_536);
  assign _zz_551 = (_zz_549 ? _zz_534 : _zz_537);
  assign _zz_552 = ((! _zz_545) || (_zz_542 && (_zz_544 <= _zz_541)));
  assign _zz_553 = (_zz_552 ? _zz_541 : _zz_544);
  assign _zz_554 = (_zz_552 ? _zz_542 : _zz_545);
  assign _zz_555 = ((! _zz_551) || (_zz_548 && (_zz_550 <= _zz_547)));
  assign _zz_556 = (_zz_555 ? _zz_547 : _zz_550);
  assign _zz_557 = (_zz_555 ? _zz_548 : _zz_551);
  assign _zz_558 = ((! _zz_557) || (_zz_554 && (_zz_556 <= _zz_553)));
  assign _zz_559 = (_zz_558 ? _zz_553 : _zz_556);
  assign _zz_560 = ((! (_zz_538 ? _zz_510 : _zz_513)) || ((_zz_558 ? _zz_554 : _zz_557) && (_zz_539 <= _zz_559)));
  assign _zz_563 = (_zz_387 < _zz_561);
  assign _zz_564 = (_zz_563 ? _zz_562 : 7'h0);
  assign io_targets = {_zz_563,{_zz_350,targets_0_iep}};
  always @ (*) begin
    io_apb_PREADY = 1'b1;
    if(_zz_708)begin
      io_apb_PREADY = 1'b0;
    end
  end

  always @ (*) begin
    io_apb_PRDATA = 32'h0;
    case(io_apb_PADDR)
      24'h0000d4 : begin
        io_apb_PRDATA[1 : 0] = gateways_0_priority;
      end
      24'h0010d4 : begin
        io_apb_PRDATA[0 : 0] = gateways_0_ip;
      end
      24'h000138 : begin
        io_apb_PRDATA[1 : 0] = gateways_1_priority;
      end
      24'h001138 : begin
        io_apb_PRDATA[0 : 0] = gateways_1_ip;
      end
      24'h00000c : begin
        io_apb_PRDATA[1 : 0] = gateways_2_priority;
      end
      24'h00100c : begin
        io_apb_PRDATA[0 : 0] = gateways_2_ip;
      end
      24'h00006c : begin
        io_apb_PRDATA[1 : 0] = gateways_3_priority;
      end
      24'h00106c : begin
        io_apb_PRDATA[0 : 0] = gateways_3_ip;
      end
      24'h0001b4 : begin
        io_apb_PRDATA[1 : 0] = gateways_4_priority;
      end
      24'h0011b4 : begin
        io_apb_PRDATA[0 : 0] = gateways_4_ip;
      end
      24'h000108 : begin
        io_apb_PRDATA[1 : 0] = gateways_5_priority;
      end
      24'h001108 : begin
        io_apb_PRDATA[0 : 0] = gateways_5_ip;
      end
      24'h000140 : begin
        io_apb_PRDATA[1 : 0] = gateways_6_priority;
      end
      24'h001140 : begin
        io_apb_PRDATA[0 : 0] = gateways_6_ip;
      end
      24'h00007c : begin
        io_apb_PRDATA[1 : 0] = gateways_7_priority;
      end
      24'h00107c : begin
        io_apb_PRDATA[0 : 0] = gateways_7_ip;
      end
      24'h0001ec : begin
        io_apb_PRDATA[1 : 0] = gateways_8_priority;
      end
      24'h0011ec : begin
        io_apb_PRDATA[0 : 0] = gateways_8_ip;
      end
      24'h0001bc : begin
        io_apb_PRDATA[1 : 0] = gateways_9_priority;
      end
      24'h0011bc : begin
        io_apb_PRDATA[0 : 0] = gateways_9_ip;
      end
      24'h000120 : begin
        io_apb_PRDATA[1 : 0] = gateways_10_priority;
      end
      24'h001120 : begin
        io_apb_PRDATA[0 : 0] = gateways_10_ip;
      end
      24'h000144 : begin
        io_apb_PRDATA[1 : 0] = gateways_11_priority;
      end
      24'h001144 : begin
        io_apb_PRDATA[0 : 0] = gateways_11_ip;
      end
      24'h000130 : begin
        io_apb_PRDATA[1 : 0] = gateways_12_priority;
      end
      24'h001130 : begin
        io_apb_PRDATA[0 : 0] = gateways_12_ip;
      end
      24'h0001b0 : begin
        io_apb_PRDATA[1 : 0] = gateways_13_priority;
      end
      24'h0011b0 : begin
        io_apb_PRDATA[0 : 0] = gateways_13_ip;
      end
      24'h0000d0 : begin
        io_apb_PRDATA[1 : 0] = gateways_14_priority;
      end
      24'h0010d0 : begin
        io_apb_PRDATA[0 : 0] = gateways_14_ip;
      end
      24'h000054 : begin
        io_apb_PRDATA[1 : 0] = gateways_15_priority;
      end
      24'h001054 : begin
        io_apb_PRDATA[0 : 0] = gateways_15_ip;
      end
      24'h000114 : begin
        io_apb_PRDATA[1 : 0] = gateways_16_priority;
      end
      24'h001114 : begin
        io_apb_PRDATA[0 : 0] = gateways_16_ip;
      end
      24'h000100 : begin
        io_apb_PRDATA[1 : 0] = gateways_17_priority;
      end
      24'h001100 : begin
        io_apb_PRDATA[0 : 0] = gateways_17_ip;
      end
      24'h0001a4 : begin
        io_apb_PRDATA[1 : 0] = gateways_18_priority;
      end
      24'h0011a4 : begin
        io_apb_PRDATA[0 : 0] = gateways_18_ip;
      end
      24'h000154 : begin
        io_apb_PRDATA[1 : 0] = gateways_19_priority;
      end
      24'h001154 : begin
        io_apb_PRDATA[0 : 0] = gateways_19_ip;
      end
      24'h00002c : begin
        io_apb_PRDATA[1 : 0] = gateways_20_priority;
      end
      24'h00102c : begin
        io_apb_PRDATA[0 : 0] = gateways_20_ip;
      end
      24'h0000e0 : begin
        io_apb_PRDATA[1 : 0] = gateways_21_priority;
      end
      24'h0010e0 : begin
        io_apb_PRDATA[0 : 0] = gateways_21_ip;
      end
      24'h000118 : begin
        io_apb_PRDATA[1 : 0] = gateways_22_priority;
      end
      24'h001118 : begin
        io_apb_PRDATA[0 : 0] = gateways_22_ip;
      end
      24'h0000c4 : begin
        io_apb_PRDATA[1 : 0] = gateways_23_priority;
      end
      24'h0010c4 : begin
        io_apb_PRDATA[0 : 0] = gateways_23_ip;
      end
      24'h000098 : begin
        io_apb_PRDATA[1 : 0] = gateways_24_priority;
      end
      24'h001098 : begin
        io_apb_PRDATA[0 : 0] = gateways_24_ip;
      end
      24'h0000fc : begin
        io_apb_PRDATA[1 : 0] = gateways_25_priority;
      end
      24'h0010fc : begin
        io_apb_PRDATA[0 : 0] = gateways_25_ip;
      end
      24'h0001a8 : begin
        io_apb_PRDATA[1 : 0] = gateways_26_priority;
      end
      24'h0011a8 : begin
        io_apb_PRDATA[0 : 0] = gateways_26_ip;
      end
      24'h000150 : begin
        io_apb_PRDATA[1 : 0] = gateways_27_priority;
      end
      24'h001150 : begin
        io_apb_PRDATA[0 : 0] = gateways_27_ip;
      end
      24'h0001c0 : begin
        io_apb_PRDATA[1 : 0] = gateways_28_priority;
      end
      24'h0011c0 : begin
        io_apb_PRDATA[0 : 0] = gateways_28_ip;
      end
      24'h000060 : begin
        io_apb_PRDATA[1 : 0] = gateways_29_priority;
      end
      24'h001060 : begin
        io_apb_PRDATA[0 : 0] = gateways_29_ip;
      end
      24'h0001f0 : begin
        io_apb_PRDATA[1 : 0] = gateways_30_priority;
      end
      24'h0011f0 : begin
        io_apb_PRDATA[0 : 0] = gateways_30_ip;
      end
      24'h000124 : begin
        io_apb_PRDATA[1 : 0] = gateways_31_priority;
      end
      24'h001124 : begin
        io_apb_PRDATA[0 : 0] = gateways_31_ip;
      end
      24'h000048 : begin
        io_apb_PRDATA[1 : 0] = gateways_32_priority;
      end
      24'h001048 : begin
        io_apb_PRDATA[0 : 0] = gateways_32_ip;
      end
      24'h00018c : begin
        io_apb_PRDATA[1 : 0] = gateways_33_priority;
      end
      24'h00118c : begin
        io_apb_PRDATA[0 : 0] = gateways_33_ip;
      end
      24'h000160 : begin
        io_apb_PRDATA[1 : 0] = gateways_34_priority;
      end
      24'h001160 : begin
        io_apb_PRDATA[0 : 0] = gateways_34_ip;
      end
      24'h200000 : begin
        io_apb_PRDATA[1 : 0] = targets_0_threshold;
      end
      24'h200004 : begin
        io_apb_PRDATA[6 : 0] = targets_0_claim;
      end
      24'h002004 : begin
        io_apb_PRDATA[21 : 21] = targets_0_ie_0;
        io_apb_PRDATA[20 : 20] = targets_0_ie_14;
        io_apb_PRDATA[24 : 24] = targets_0_ie_21;
        io_apb_PRDATA[17 : 17] = targets_0_ie_23;
        io_apb_PRDATA[6 : 6] = targets_0_ie_24;
        io_apb_PRDATA[31 : 31] = targets_0_ie_25;
      end
      24'h002008 : begin
        io_apb_PRDATA[14 : 14] = targets_0_ie_1;
        io_apb_PRDATA[2 : 2] = targets_0_ie_5;
        io_apb_PRDATA[16 : 16] = targets_0_ie_6;
        io_apb_PRDATA[8 : 8] = targets_0_ie_10;
        io_apb_PRDATA[17 : 17] = targets_0_ie_11;
        io_apb_PRDATA[12 : 12] = targets_0_ie_12;
        io_apb_PRDATA[5 : 5] = targets_0_ie_16;
        io_apb_PRDATA[0 : 0] = targets_0_ie_17;
        io_apb_PRDATA[21 : 21] = targets_0_ie_19;
        io_apb_PRDATA[6 : 6] = targets_0_ie_22;
        io_apb_PRDATA[20 : 20] = targets_0_ie_27;
        io_apb_PRDATA[9 : 9] = targets_0_ie_31;
        io_apb_PRDATA[24 : 24] = targets_0_ie_34;
      end
      24'h002000 : begin
        io_apb_PRDATA[3 : 3] = targets_0_ie_2;
        io_apb_PRDATA[27 : 27] = targets_0_ie_3;
        io_apb_PRDATA[31 : 31] = targets_0_ie_7;
        io_apb_PRDATA[21 : 21] = targets_0_ie_15;
        io_apb_PRDATA[11 : 11] = targets_0_ie_20;
        io_apb_PRDATA[24 : 24] = targets_0_ie_29;
        io_apb_PRDATA[18 : 18] = targets_0_ie_32;
      end
      24'h00200c : begin
        io_apb_PRDATA[13 : 13] = targets_0_ie_4;
        io_apb_PRDATA[27 : 27] = targets_0_ie_8;
        io_apb_PRDATA[15 : 15] = targets_0_ie_9;
        io_apb_PRDATA[12 : 12] = targets_0_ie_13;
        io_apb_PRDATA[9 : 9] = targets_0_ie_18;
        io_apb_PRDATA[10 : 10] = targets_0_ie_26;
        io_apb_PRDATA[16 : 16] = targets_0_ie_28;
        io_apb_PRDATA[28 : 28] = targets_0_ie_30;
        io_apb_PRDATA[3 : 3] = targets_0_ie_33;
      end
      24'h201000 : begin
        io_apb_PRDATA[1 : 0] = _zz_174;
      end
      24'h201004 : begin
        io_apb_PRDATA[6 : 0] = _zz_351;
      end
      24'h002084 : begin
        io_apb_PRDATA[21 : 21] = _zz_139;
        io_apb_PRDATA[20 : 20] = _zz_153;
        io_apb_PRDATA[24 : 24] = _zz_160;
        io_apb_PRDATA[17 : 17] = _zz_162;
        io_apb_PRDATA[6 : 6] = _zz_163;
        io_apb_PRDATA[31 : 31] = _zz_164;
      end
      24'h002088 : begin
        io_apb_PRDATA[14 : 14] = _zz_140;
        io_apb_PRDATA[2 : 2] = _zz_144;
        io_apb_PRDATA[16 : 16] = _zz_145;
        io_apb_PRDATA[8 : 8] = _zz_149;
        io_apb_PRDATA[17 : 17] = _zz_150;
        io_apb_PRDATA[12 : 12] = _zz_151;
        io_apb_PRDATA[5 : 5] = _zz_155;
        io_apb_PRDATA[0 : 0] = _zz_156;
        io_apb_PRDATA[21 : 21] = _zz_158;
        io_apb_PRDATA[6 : 6] = _zz_161;
        io_apb_PRDATA[20 : 20] = _zz_166;
        io_apb_PRDATA[9 : 9] = _zz_170;
        io_apb_PRDATA[24 : 24] = _zz_173;
      end
      24'h002080 : begin
        io_apb_PRDATA[3 : 3] = _zz_141;
        io_apb_PRDATA[27 : 27] = _zz_142;
        io_apb_PRDATA[31 : 31] = _zz_146;
        io_apb_PRDATA[21 : 21] = _zz_154;
        io_apb_PRDATA[11 : 11] = _zz_159;
        io_apb_PRDATA[24 : 24] = _zz_168;
        io_apb_PRDATA[18 : 18] = _zz_171;
      end
      24'h00208c : begin
        io_apb_PRDATA[13 : 13] = _zz_143;
        io_apb_PRDATA[27 : 27] = _zz_147;
        io_apb_PRDATA[15 : 15] = _zz_148;
        io_apb_PRDATA[12 : 12] = _zz_152;
        io_apb_PRDATA[9 : 9] = _zz_157;
        io_apb_PRDATA[10 : 10] = _zz_165;
        io_apb_PRDATA[16 : 16] = _zz_167;
        io_apb_PRDATA[28 : 28] = _zz_169;
        io_apb_PRDATA[3 : 3] = _zz_172;
      end
      24'h202000 : begin
        io_apb_PRDATA[1 : 0] = _zz_387;
      end
      24'h202004 : begin
        io_apb_PRDATA[6 : 0] = _zz_564;
      end
      24'h002104 : begin
        io_apb_PRDATA[21 : 21] = _zz_352;
        io_apb_PRDATA[20 : 20] = _zz_366;
        io_apb_PRDATA[24 : 24] = _zz_373;
        io_apb_PRDATA[17 : 17] = _zz_375;
        io_apb_PRDATA[6 : 6] = _zz_376;
        io_apb_PRDATA[31 : 31] = _zz_377;
      end
      24'h002108 : begin
        io_apb_PRDATA[14 : 14] = _zz_353;
        io_apb_PRDATA[2 : 2] = _zz_357;
        io_apb_PRDATA[16 : 16] = _zz_358;
        io_apb_PRDATA[8 : 8] = _zz_362;
        io_apb_PRDATA[17 : 17] = _zz_363;
        io_apb_PRDATA[12 : 12] = _zz_364;
        io_apb_PRDATA[5 : 5] = _zz_368;
        io_apb_PRDATA[0 : 0] = _zz_369;
        io_apb_PRDATA[21 : 21] = _zz_371;
        io_apb_PRDATA[6 : 6] = _zz_374;
        io_apb_PRDATA[20 : 20] = _zz_379;
        io_apb_PRDATA[9 : 9] = _zz_383;
        io_apb_PRDATA[24 : 24] = _zz_386;
      end
      24'h002100 : begin
        io_apb_PRDATA[3 : 3] = _zz_354;
        io_apb_PRDATA[27 : 27] = _zz_355;
        io_apb_PRDATA[31 : 31] = _zz_359;
        io_apb_PRDATA[21 : 21] = _zz_367;
        io_apb_PRDATA[11 : 11] = _zz_372;
        io_apb_PRDATA[24 : 24] = _zz_381;
        io_apb_PRDATA[18 : 18] = _zz_384;
      end
      24'h00210c : begin
        io_apb_PRDATA[13 : 13] = _zz_356;
        io_apb_PRDATA[27 : 27] = _zz_360;
        io_apb_PRDATA[15 : 15] = _zz_361;
        io_apb_PRDATA[12 : 12] = _zz_365;
        io_apb_PRDATA[9 : 9] = _zz_370;
        io_apb_PRDATA[10 : 10] = _zz_378;
        io_apb_PRDATA[16 : 16] = _zz_380;
        io_apb_PRDATA[28 : 28] = _zz_382;
        io_apb_PRDATA[3 : 3] = _zz_385;
      end
      default : begin
      end
    endcase
  end

  assign io_apb_PSLVERROR = 1'b0;
  assign bus_askWrite = ((io_apb_PSEL[0] && io_apb_PENABLE) && io_apb_PWRITE);
  assign bus_askRead = ((io_apb_PSEL[0] && io_apb_PENABLE) && (! io_apb_PWRITE));
  assign bus_doWrite = (((io_apb_PSEL[0] && io_apb_PENABLE) && io_apb_PREADY) && io_apb_PWRITE);
  assign bus_doRead = (((io_apb_PSEL[0] && io_apb_PENABLE) && io_apb_PREADY) && (! io_apb_PWRITE));
  assign gateways_0_priority = _zz_565;
  assign gateways_1_priority = _zz_566;
  assign gateways_2_priority = _zz_567;
  assign gateways_3_priority = _zz_568;
  assign gateways_4_priority = _zz_569;
  assign gateways_5_priority = _zz_570;
  assign gateways_6_priority = _zz_571;
  assign gateways_7_priority = _zz_572;
  assign gateways_8_priority = _zz_573;
  assign gateways_9_priority = _zz_574;
  assign gateways_10_priority = _zz_575;
  assign gateways_11_priority = _zz_576;
  assign gateways_12_priority = _zz_577;
  assign gateways_13_priority = _zz_578;
  assign gateways_14_priority = _zz_579;
  assign gateways_15_priority = _zz_580;
  assign gateways_16_priority = _zz_581;
  assign gateways_17_priority = _zz_582;
  assign gateways_18_priority = _zz_583;
  assign gateways_19_priority = _zz_584;
  assign gateways_20_priority = _zz_585;
  assign gateways_21_priority = _zz_586;
  assign gateways_22_priority = _zz_587;
  assign gateways_23_priority = _zz_588;
  assign gateways_24_priority = _zz_589;
  assign gateways_25_priority = _zz_590;
  assign gateways_26_priority = _zz_591;
  assign gateways_27_priority = _zz_592;
  assign gateways_28_priority = _zz_593;
  assign gateways_29_priority = _zz_594;
  assign gateways_30_priority = _zz_595;
  assign gateways_31_priority = _zz_596;
  assign gateways_32_priority = _zz_597;
  assign gateways_33_priority = _zz_598;
  assign gateways_34_priority = _zz_599;
  always @ (*) begin
    mapping_claim_valid = 1'b0;
    case(io_apb_PADDR)
      24'h200004 : begin
        if(bus_doRead)begin
          mapping_claim_valid = 1'b1;
        end
      end
      24'h201004 : begin
        if(bus_doRead)begin
          mapping_claim_valid = 1'b1;
        end
      end
      24'h202004 : begin
        if(bus_doRead)begin
          mapping_claim_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @ (*) begin
    mapping_claim_payload = 7'h0;
    case(io_apb_PADDR)
      24'h200004 : begin
        if(bus_doRead)begin
          mapping_claim_payload = targets_0_claim;
        end
      end
      24'h201004 : begin
        if(bus_doRead)begin
          mapping_claim_payload = _zz_351;
        end
      end
      24'h202004 : begin
        if(bus_doRead)begin
          mapping_claim_payload = _zz_564;
        end
      end
      default : begin
      end
    endcase
  end

  always @ (*) begin
    mapping_completion_valid = 1'b0;
    if(mapping_targetMapping_0_targetCompletion_valid)begin
      mapping_completion_valid = 1'b1;
    end
    if(mapping_targetMapping_1_targetCompletion_valid)begin
      mapping_completion_valid = 1'b1;
    end
    if(mapping_targetMapping_2_targetCompletion_valid)begin
      mapping_completion_valid = 1'b1;
    end
  end

  always @ (*) begin
    mapping_completion_payload = 7'h0;
    if(mapping_targetMapping_0_targetCompletion_valid)begin
      mapping_completion_payload = mapping_targetMapping_0_targetCompletion_payload;
    end
    if(mapping_targetMapping_1_targetCompletion_valid)begin
      mapping_completion_payload = mapping_targetMapping_1_targetCompletion_payload;
    end
    if(mapping_targetMapping_2_targetCompletion_valid)begin
      mapping_completion_payload = mapping_targetMapping_2_targetCompletion_payload;
    end
  end

  always @ (*) begin
    mapping_coherencyStall_willIncrement = 1'b0;
    if(_zz_708)begin
      mapping_coherencyStall_willIncrement = 1'b1;
    end
    if(1'b1)begin
      if(bus_askWrite)begin
        mapping_coherencyStall_willIncrement = 1'b1;
      end
      if(bus_askRead)begin
        mapping_coherencyStall_willIncrement = 1'b1;
      end
    end
  end

  assign mapping_coherencyStall_willClear = 1'b0;
  assign mapping_coherencyStall_willOverflowIfInc = (mapping_coherencyStall_value == 1'b1);
  assign mapping_coherencyStall_willOverflow = (mapping_coherencyStall_willOverflowIfInc && mapping_coherencyStall_willIncrement);
  always @ (*) begin
    mapping_coherencyStall_valueNext = (mapping_coherencyStall_value + mapping_coherencyStall_willIncrement);
    if(mapping_coherencyStall_willClear)begin
      mapping_coherencyStall_valueNext = 1'b0;
    end
  end

  assign targets_0_threshold = _zz_600;
  always @ (*) begin
    mapping_targetMapping_0_targetCompletion_valid = 1'b0;
    case(io_apb_PADDR)
      24'h200004 : begin
        if(bus_doWrite)begin
          mapping_targetMapping_0_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign targets_0_ie_0 = _zz_601;
  assign targets_0_ie_1 = _zz_602;
  assign targets_0_ie_2 = _zz_603;
  assign targets_0_ie_3 = _zz_604;
  assign targets_0_ie_4 = _zz_605;
  assign targets_0_ie_5 = _zz_606;
  assign targets_0_ie_6 = _zz_607;
  assign targets_0_ie_7 = _zz_608;
  assign targets_0_ie_8 = _zz_609;
  assign targets_0_ie_9 = _zz_610;
  assign targets_0_ie_10 = _zz_611;
  assign targets_0_ie_11 = _zz_612;
  assign targets_0_ie_12 = _zz_613;
  assign targets_0_ie_13 = _zz_614;
  assign targets_0_ie_14 = _zz_615;
  assign targets_0_ie_15 = _zz_616;
  assign targets_0_ie_16 = _zz_617;
  assign targets_0_ie_17 = _zz_618;
  assign targets_0_ie_18 = _zz_619;
  assign targets_0_ie_19 = _zz_620;
  assign targets_0_ie_20 = _zz_621;
  assign targets_0_ie_21 = _zz_622;
  assign targets_0_ie_22 = _zz_623;
  assign targets_0_ie_23 = _zz_624;
  assign targets_0_ie_24 = _zz_625;
  assign targets_0_ie_25 = _zz_626;
  assign targets_0_ie_26 = _zz_627;
  assign targets_0_ie_27 = _zz_628;
  assign targets_0_ie_28 = _zz_629;
  assign targets_0_ie_29 = _zz_630;
  assign targets_0_ie_30 = _zz_631;
  assign targets_0_ie_31 = _zz_632;
  assign targets_0_ie_32 = _zz_633;
  assign targets_0_ie_33 = _zz_634;
  assign targets_0_ie_34 = _zz_635;
  assign _zz_174 = _zz_636;
  always @ (*) begin
    mapping_targetMapping_1_targetCompletion_valid = 1'b0;
    case(io_apb_PADDR)
      24'h201004 : begin
        if(bus_doWrite)begin
          mapping_targetMapping_1_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign _zz_139 = _zz_637;
  assign _zz_140 = _zz_638;
  assign _zz_141 = _zz_639;
  assign _zz_142 = _zz_640;
  assign _zz_143 = _zz_641;
  assign _zz_144 = _zz_642;
  assign _zz_145 = _zz_643;
  assign _zz_146 = _zz_644;
  assign _zz_147 = _zz_645;
  assign _zz_148 = _zz_646;
  assign _zz_149 = _zz_647;
  assign _zz_150 = _zz_648;
  assign _zz_151 = _zz_649;
  assign _zz_152 = _zz_650;
  assign _zz_153 = _zz_651;
  assign _zz_154 = _zz_652;
  assign _zz_155 = _zz_653;
  assign _zz_156 = _zz_654;
  assign _zz_157 = _zz_655;
  assign _zz_158 = _zz_656;
  assign _zz_159 = _zz_657;
  assign _zz_160 = _zz_658;
  assign _zz_161 = _zz_659;
  assign _zz_162 = _zz_660;
  assign _zz_163 = _zz_661;
  assign _zz_164 = _zz_662;
  assign _zz_165 = _zz_663;
  assign _zz_166 = _zz_664;
  assign _zz_167 = _zz_665;
  assign _zz_168 = _zz_666;
  assign _zz_169 = _zz_667;
  assign _zz_170 = _zz_668;
  assign _zz_171 = _zz_669;
  assign _zz_172 = _zz_670;
  assign _zz_173 = _zz_671;
  assign _zz_387 = _zz_672;
  always @ (*) begin
    mapping_targetMapping_2_targetCompletion_valid = 1'b0;
    case(io_apb_PADDR)
      24'h202004 : begin
        if(bus_doWrite)begin
          mapping_targetMapping_2_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign _zz_352 = _zz_673;
  assign _zz_353 = _zz_674;
  assign _zz_354 = _zz_675;
  assign _zz_355 = _zz_676;
  assign _zz_356 = _zz_677;
  assign _zz_357 = _zz_678;
  assign _zz_358 = _zz_679;
  assign _zz_359 = _zz_680;
  assign _zz_360 = _zz_681;
  assign _zz_361 = _zz_682;
  assign _zz_362 = _zz_683;
  assign _zz_363 = _zz_684;
  assign _zz_364 = _zz_685;
  assign _zz_365 = _zz_686;
  assign _zz_366 = _zz_687;
  assign _zz_367 = _zz_688;
  assign _zz_368 = _zz_689;
  assign _zz_369 = _zz_690;
  assign _zz_370 = _zz_691;
  assign _zz_371 = _zz_692;
  assign _zz_372 = _zz_693;
  assign _zz_373 = _zz_694;
  assign _zz_374 = _zz_695;
  assign _zz_375 = _zz_696;
  assign _zz_376 = _zz_697;
  assign _zz_377 = _zz_698;
  assign _zz_378 = _zz_699;
  assign _zz_379 = _zz_700;
  assign _zz_380 = _zz_701;
  assign _zz_381 = _zz_702;
  assign _zz_382 = _zz_703;
  assign _zz_383 = _zz_704;
  assign _zz_384 = _zz_705;
  assign _zz_385 = _zz_706;
  assign _zz_386 = _zz_707;
  assign mapping_targetMapping_0_targetCompletion_payload = io_apb_PWDATA[6 : 0];
  assign mapping_targetMapping_1_targetCompletion_payload = io_apb_PWDATA[6 : 0];
  assign mapping_targetMapping_2_targetCompletion_payload = io_apb_PWDATA[6 : 0];
  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      gateways_0_ip <= 1'b0;
      gateways_0_waitCompletion <= 1'b0;
      gateways_1_ip <= 1'b0;
      gateways_1_waitCompletion <= 1'b0;
      gateways_2_ip <= 1'b0;
      gateways_2_waitCompletion <= 1'b0;
      gateways_3_ip <= 1'b0;
      gateways_3_waitCompletion <= 1'b0;
      gateways_4_ip <= 1'b0;
      gateways_4_waitCompletion <= 1'b0;
      gateways_5_ip <= 1'b0;
      gateways_5_waitCompletion <= 1'b0;
      gateways_6_ip <= 1'b0;
      gateways_6_waitCompletion <= 1'b0;
      gateways_7_ip <= 1'b0;
      gateways_7_waitCompletion <= 1'b0;
      gateways_8_ip <= 1'b0;
      gateways_8_waitCompletion <= 1'b0;
      gateways_9_ip <= 1'b0;
      gateways_9_waitCompletion <= 1'b0;
      gateways_10_ip <= 1'b0;
      gateways_10_waitCompletion <= 1'b0;
      gateways_11_ip <= 1'b0;
      gateways_11_waitCompletion <= 1'b0;
      gateways_12_ip <= 1'b0;
      gateways_12_waitCompletion <= 1'b0;
      gateways_13_ip <= 1'b0;
      gateways_13_waitCompletion <= 1'b0;
      gateways_14_ip <= 1'b0;
      gateways_14_waitCompletion <= 1'b0;
      gateways_15_ip <= 1'b0;
      gateways_15_waitCompletion <= 1'b0;
      gateways_16_ip <= 1'b0;
      gateways_16_waitCompletion <= 1'b0;
      gateways_17_ip <= 1'b0;
      gateways_17_waitCompletion <= 1'b0;
      gateways_18_ip <= 1'b0;
      gateways_18_waitCompletion <= 1'b0;
      gateways_19_ip <= 1'b0;
      gateways_19_waitCompletion <= 1'b0;
      gateways_20_ip <= 1'b0;
      gateways_20_waitCompletion <= 1'b0;
      gateways_21_ip <= 1'b0;
      gateways_21_waitCompletion <= 1'b0;
      gateways_22_ip <= 1'b0;
      gateways_22_waitCompletion <= 1'b0;
      gateways_23_ip <= 1'b0;
      gateways_23_waitCompletion <= 1'b0;
      gateways_24_ip <= 1'b0;
      gateways_24_waitCompletion <= 1'b0;
      gateways_25_ip <= 1'b0;
      gateways_25_waitCompletion <= 1'b0;
      gateways_26_ip <= 1'b0;
      gateways_26_waitCompletion <= 1'b0;
      gateways_27_ip <= 1'b0;
      gateways_27_waitCompletion <= 1'b0;
      gateways_28_ip <= 1'b0;
      gateways_28_waitCompletion <= 1'b0;
      gateways_29_ip <= 1'b0;
      gateways_29_waitCompletion <= 1'b0;
      gateways_30_ip <= 1'b0;
      gateways_30_waitCompletion <= 1'b0;
      gateways_31_ip <= 1'b0;
      gateways_31_waitCompletion <= 1'b0;
      gateways_32_ip <= 1'b0;
      gateways_32_waitCompletion <= 1'b0;
      gateways_33_ip <= 1'b0;
      gateways_33_waitCompletion <= 1'b0;
      gateways_34_ip <= 1'b0;
      gateways_34_waitCompletion <= 1'b0;
      _zz_565 <= 2'b00;
      _zz_566 <= 2'b00;
      _zz_567 <= 2'b00;
      _zz_568 <= 2'b00;
      _zz_569 <= 2'b00;
      _zz_570 <= 2'b00;
      _zz_571 <= 2'b00;
      _zz_572 <= 2'b00;
      _zz_573 <= 2'b00;
      _zz_574 <= 2'b00;
      _zz_575 <= 2'b00;
      _zz_576 <= 2'b00;
      _zz_577 <= 2'b00;
      _zz_578 <= 2'b00;
      _zz_579 <= 2'b00;
      _zz_580 <= 2'b00;
      _zz_581 <= 2'b00;
      _zz_582 <= 2'b00;
      _zz_583 <= 2'b00;
      _zz_584 <= 2'b00;
      _zz_585 <= 2'b00;
      _zz_586 <= 2'b00;
      _zz_587 <= 2'b00;
      _zz_588 <= 2'b00;
      _zz_589 <= 2'b00;
      _zz_590 <= 2'b00;
      _zz_591 <= 2'b00;
      _zz_592 <= 2'b00;
      _zz_593 <= 2'b00;
      _zz_594 <= 2'b00;
      _zz_595 <= 2'b00;
      _zz_596 <= 2'b00;
      _zz_597 <= 2'b00;
      _zz_598 <= 2'b00;
      _zz_599 <= 2'b00;
      mapping_coherencyStall_value <= 1'b0;
      _zz_600 <= 2'b00;
      _zz_601 <= 1'b0;
      _zz_602 <= 1'b0;
      _zz_603 <= 1'b0;
      _zz_604 <= 1'b0;
      _zz_605 <= 1'b0;
      _zz_606 <= 1'b0;
      _zz_607 <= 1'b0;
      _zz_608 <= 1'b0;
      _zz_609 <= 1'b0;
      _zz_610 <= 1'b0;
      _zz_611 <= 1'b0;
      _zz_612 <= 1'b0;
      _zz_613 <= 1'b0;
      _zz_614 <= 1'b0;
      _zz_615 <= 1'b0;
      _zz_616 <= 1'b0;
      _zz_617 <= 1'b0;
      _zz_618 <= 1'b0;
      _zz_619 <= 1'b0;
      _zz_620 <= 1'b0;
      _zz_621 <= 1'b0;
      _zz_622 <= 1'b0;
      _zz_623 <= 1'b0;
      _zz_624 <= 1'b0;
      _zz_625 <= 1'b0;
      _zz_626 <= 1'b0;
      _zz_627 <= 1'b0;
      _zz_628 <= 1'b0;
      _zz_629 <= 1'b0;
      _zz_630 <= 1'b0;
      _zz_631 <= 1'b0;
      _zz_632 <= 1'b0;
      _zz_633 <= 1'b0;
      _zz_634 <= 1'b0;
      _zz_635 <= 1'b0;
      _zz_636 <= 2'b00;
      _zz_637 <= 1'b0;
      _zz_638 <= 1'b0;
      _zz_639 <= 1'b0;
      _zz_640 <= 1'b0;
      _zz_641 <= 1'b0;
      _zz_642 <= 1'b0;
      _zz_643 <= 1'b0;
      _zz_644 <= 1'b0;
      _zz_645 <= 1'b0;
      _zz_646 <= 1'b0;
      _zz_647 <= 1'b0;
      _zz_648 <= 1'b0;
      _zz_649 <= 1'b0;
      _zz_650 <= 1'b0;
      _zz_651 <= 1'b0;
      _zz_652 <= 1'b0;
      _zz_653 <= 1'b0;
      _zz_654 <= 1'b0;
      _zz_655 <= 1'b0;
      _zz_656 <= 1'b0;
      _zz_657 <= 1'b0;
      _zz_658 <= 1'b0;
      _zz_659 <= 1'b0;
      _zz_660 <= 1'b0;
      _zz_661 <= 1'b0;
      _zz_662 <= 1'b0;
      _zz_663 <= 1'b0;
      _zz_664 <= 1'b0;
      _zz_665 <= 1'b0;
      _zz_666 <= 1'b0;
      _zz_667 <= 1'b0;
      _zz_668 <= 1'b0;
      _zz_669 <= 1'b0;
      _zz_670 <= 1'b0;
      _zz_671 <= 1'b0;
      _zz_672 <= 2'b00;
      _zz_673 <= 1'b0;
      _zz_674 <= 1'b0;
      _zz_675 <= 1'b0;
      _zz_676 <= 1'b0;
      _zz_677 <= 1'b0;
      _zz_678 <= 1'b0;
      _zz_679 <= 1'b0;
      _zz_680 <= 1'b0;
      _zz_681 <= 1'b0;
      _zz_682 <= 1'b0;
      _zz_683 <= 1'b0;
      _zz_684 <= 1'b0;
      _zz_685 <= 1'b0;
      _zz_686 <= 1'b0;
      _zz_687 <= 1'b0;
      _zz_688 <= 1'b0;
      _zz_689 <= 1'b0;
      _zz_690 <= 1'b0;
      _zz_691 <= 1'b0;
      _zz_692 <= 1'b0;
      _zz_693 <= 1'b0;
      _zz_694 <= 1'b0;
      _zz_695 <= 1'b0;
      _zz_696 <= 1'b0;
      _zz_697 <= 1'b0;
      _zz_698 <= 1'b0;
      _zz_699 <= 1'b0;
      _zz_700 <= 1'b0;
      _zz_701 <= 1'b0;
      _zz_702 <= 1'b0;
      _zz_703 <= 1'b0;
      _zz_704 <= 1'b0;
      _zz_705 <= 1'b0;
      _zz_706 <= 1'b0;
      _zz_707 <= 1'b0;
    end else begin
      if((! gateways_0_waitCompletion))begin
        gateways_0_ip <= _zz_1;
        gateways_0_waitCompletion <= _zz_1;
      end
      if((! gateways_1_waitCompletion))begin
        gateways_1_ip <= _zz_2;
        gateways_1_waitCompletion <= _zz_2;
      end
      if((! gateways_2_waitCompletion))begin
        gateways_2_ip <= _zz_3;
        gateways_2_waitCompletion <= _zz_3;
      end
      if((! gateways_3_waitCompletion))begin
        gateways_3_ip <= _zz_4;
        gateways_3_waitCompletion <= _zz_4;
      end
      if((! gateways_4_waitCompletion))begin
        gateways_4_ip <= _zz_5;
        gateways_4_waitCompletion <= _zz_5;
      end
      if((! gateways_5_waitCompletion))begin
        gateways_5_ip <= _zz_6;
        gateways_5_waitCompletion <= _zz_6;
      end
      if((! gateways_6_waitCompletion))begin
        gateways_6_ip <= _zz_7;
        gateways_6_waitCompletion <= _zz_7;
      end
      if((! gateways_7_waitCompletion))begin
        gateways_7_ip <= _zz_8;
        gateways_7_waitCompletion <= _zz_8;
      end
      if((! gateways_8_waitCompletion))begin
        gateways_8_ip <= _zz_9;
        gateways_8_waitCompletion <= _zz_9;
      end
      if((! gateways_9_waitCompletion))begin
        gateways_9_ip <= _zz_10;
        gateways_9_waitCompletion <= _zz_10;
      end
      if((! gateways_10_waitCompletion))begin
        gateways_10_ip <= _zz_11;
        gateways_10_waitCompletion <= _zz_11;
      end
      if((! gateways_11_waitCompletion))begin
        gateways_11_ip <= _zz_12;
        gateways_11_waitCompletion <= _zz_12;
      end
      if((! gateways_12_waitCompletion))begin
        gateways_12_ip <= _zz_13;
        gateways_12_waitCompletion <= _zz_13;
      end
      if((! gateways_13_waitCompletion))begin
        gateways_13_ip <= _zz_14;
        gateways_13_waitCompletion <= _zz_14;
      end
      if((! gateways_14_waitCompletion))begin
        gateways_14_ip <= _zz_15;
        gateways_14_waitCompletion <= _zz_15;
      end
      if((! gateways_15_waitCompletion))begin
        gateways_15_ip <= _zz_16;
        gateways_15_waitCompletion <= _zz_16;
      end
      if((! gateways_16_waitCompletion))begin
        gateways_16_ip <= _zz_17;
        gateways_16_waitCompletion <= _zz_17;
      end
      if((! gateways_17_waitCompletion))begin
        gateways_17_ip <= _zz_18;
        gateways_17_waitCompletion <= _zz_18;
      end
      if((! gateways_18_waitCompletion))begin
        gateways_18_ip <= _zz_19;
        gateways_18_waitCompletion <= _zz_19;
      end
      if((! gateways_19_waitCompletion))begin
        gateways_19_ip <= _zz_20;
        gateways_19_waitCompletion <= _zz_20;
      end
      if((! gateways_20_waitCompletion))begin
        gateways_20_ip <= _zz_21;
        gateways_20_waitCompletion <= _zz_21;
      end
      if((! gateways_21_waitCompletion))begin
        gateways_21_ip <= _zz_22;
        gateways_21_waitCompletion <= _zz_22;
      end
      if((! gateways_22_waitCompletion))begin
        gateways_22_ip <= _zz_23;
        gateways_22_waitCompletion <= _zz_23;
      end
      if((! gateways_23_waitCompletion))begin
        gateways_23_ip <= _zz_24;
        gateways_23_waitCompletion <= _zz_24;
      end
      if((! gateways_24_waitCompletion))begin
        gateways_24_ip <= _zz_25;
        gateways_24_waitCompletion <= _zz_25;
      end
      if((! gateways_25_waitCompletion))begin
        gateways_25_ip <= _zz_26;
        gateways_25_waitCompletion <= _zz_26;
      end
      if((! gateways_26_waitCompletion))begin
        gateways_26_ip <= _zz_27;
        gateways_26_waitCompletion <= _zz_27;
      end
      if((! gateways_27_waitCompletion))begin
        gateways_27_ip <= _zz_28;
        gateways_27_waitCompletion <= _zz_28;
      end
      if((! gateways_28_waitCompletion))begin
        gateways_28_ip <= _zz_29;
        gateways_28_waitCompletion <= _zz_29;
      end
      if((! gateways_29_waitCompletion))begin
        gateways_29_ip <= _zz_30;
        gateways_29_waitCompletion <= _zz_30;
      end
      if((! gateways_30_waitCompletion))begin
        gateways_30_ip <= _zz_31;
        gateways_30_waitCompletion <= _zz_31;
      end
      if((! gateways_31_waitCompletion))begin
        gateways_31_ip <= _zz_32;
        gateways_31_waitCompletion <= _zz_32;
      end
      if((! gateways_32_waitCompletion))begin
        gateways_32_ip <= _zz_33;
        gateways_32_waitCompletion <= _zz_33;
      end
      if((! gateways_33_waitCompletion))begin
        gateways_33_ip <= _zz_34;
        gateways_33_waitCompletion <= _zz_34;
      end
      if((! gateways_34_waitCompletion))begin
        gateways_34_ip <= _zz_35;
        gateways_34_waitCompletion <= _zz_35;
      end
      if(mapping_claim_valid)begin
        case(mapping_claim_payload)
          7'h35 : begin
            gateways_0_ip <= 1'b0;
          end
          7'h4e : begin
            gateways_1_ip <= 1'b0;
          end
          7'h03 : begin
            gateways_2_ip <= 1'b0;
          end
          7'h1b : begin
            gateways_3_ip <= 1'b0;
          end
          7'h6d : begin
            gateways_4_ip <= 1'b0;
          end
          7'h42 : begin
            gateways_5_ip <= 1'b0;
          end
          7'h50 : begin
            gateways_6_ip <= 1'b0;
          end
          7'h1f : begin
            gateways_7_ip <= 1'b0;
          end
          7'h7b : begin
            gateways_8_ip <= 1'b0;
          end
          7'h6f : begin
            gateways_9_ip <= 1'b0;
          end
          7'h48 : begin
            gateways_10_ip <= 1'b0;
          end
          7'h51 : begin
            gateways_11_ip <= 1'b0;
          end
          7'h4c : begin
            gateways_12_ip <= 1'b0;
          end
          7'h6c : begin
            gateways_13_ip <= 1'b0;
          end
          7'h34 : begin
            gateways_14_ip <= 1'b0;
          end
          7'h15 : begin
            gateways_15_ip <= 1'b0;
          end
          7'h45 : begin
            gateways_16_ip <= 1'b0;
          end
          7'h40 : begin
            gateways_17_ip <= 1'b0;
          end
          7'h69 : begin
            gateways_18_ip <= 1'b0;
          end
          7'h55 : begin
            gateways_19_ip <= 1'b0;
          end
          7'h0b : begin
            gateways_20_ip <= 1'b0;
          end
          7'h38 : begin
            gateways_21_ip <= 1'b0;
          end
          7'h46 : begin
            gateways_22_ip <= 1'b0;
          end
          7'h31 : begin
            gateways_23_ip <= 1'b0;
          end
          7'h26 : begin
            gateways_24_ip <= 1'b0;
          end
          7'h3f : begin
            gateways_25_ip <= 1'b0;
          end
          7'h6a : begin
            gateways_26_ip <= 1'b0;
          end
          7'h54 : begin
            gateways_27_ip <= 1'b0;
          end
          7'h70 : begin
            gateways_28_ip <= 1'b0;
          end
          7'h18 : begin
            gateways_29_ip <= 1'b0;
          end
          7'h7c : begin
            gateways_30_ip <= 1'b0;
          end
          7'h49 : begin
            gateways_31_ip <= 1'b0;
          end
          7'h12 : begin
            gateways_32_ip <= 1'b0;
          end
          7'h63 : begin
            gateways_33_ip <= 1'b0;
          end
          7'h58 : begin
            gateways_34_ip <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      if(mapping_completion_valid)begin
        case(mapping_completion_payload)
          7'h35 : begin
            gateways_0_waitCompletion <= 1'b0;
          end
          7'h4e : begin
            gateways_1_waitCompletion <= 1'b0;
          end
          7'h03 : begin
            gateways_2_waitCompletion <= 1'b0;
          end
          7'h1b : begin
            gateways_3_waitCompletion <= 1'b0;
          end
          7'h6d : begin
            gateways_4_waitCompletion <= 1'b0;
          end
          7'h42 : begin
            gateways_5_waitCompletion <= 1'b0;
          end
          7'h50 : begin
            gateways_6_waitCompletion <= 1'b0;
          end
          7'h1f : begin
            gateways_7_waitCompletion <= 1'b0;
          end
          7'h7b : begin
            gateways_8_waitCompletion <= 1'b0;
          end
          7'h6f : begin
            gateways_9_waitCompletion <= 1'b0;
          end
          7'h48 : begin
            gateways_10_waitCompletion <= 1'b0;
          end
          7'h51 : begin
            gateways_11_waitCompletion <= 1'b0;
          end
          7'h4c : begin
            gateways_12_waitCompletion <= 1'b0;
          end
          7'h6c : begin
            gateways_13_waitCompletion <= 1'b0;
          end
          7'h34 : begin
            gateways_14_waitCompletion <= 1'b0;
          end
          7'h15 : begin
            gateways_15_waitCompletion <= 1'b0;
          end
          7'h45 : begin
            gateways_16_waitCompletion <= 1'b0;
          end
          7'h40 : begin
            gateways_17_waitCompletion <= 1'b0;
          end
          7'h69 : begin
            gateways_18_waitCompletion <= 1'b0;
          end
          7'h55 : begin
            gateways_19_waitCompletion <= 1'b0;
          end
          7'h0b : begin
            gateways_20_waitCompletion <= 1'b0;
          end
          7'h38 : begin
            gateways_21_waitCompletion <= 1'b0;
          end
          7'h46 : begin
            gateways_22_waitCompletion <= 1'b0;
          end
          7'h31 : begin
            gateways_23_waitCompletion <= 1'b0;
          end
          7'h26 : begin
            gateways_24_waitCompletion <= 1'b0;
          end
          7'h3f : begin
            gateways_25_waitCompletion <= 1'b0;
          end
          7'h6a : begin
            gateways_26_waitCompletion <= 1'b0;
          end
          7'h54 : begin
            gateways_27_waitCompletion <= 1'b0;
          end
          7'h70 : begin
            gateways_28_waitCompletion <= 1'b0;
          end
          7'h18 : begin
            gateways_29_waitCompletion <= 1'b0;
          end
          7'h7c : begin
            gateways_30_waitCompletion <= 1'b0;
          end
          7'h49 : begin
            gateways_31_waitCompletion <= 1'b0;
          end
          7'h12 : begin
            gateways_32_waitCompletion <= 1'b0;
          end
          7'h63 : begin
            gateways_33_waitCompletion <= 1'b0;
          end
          7'h58 : begin
            gateways_34_waitCompletion <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      mapping_coherencyStall_value <= mapping_coherencyStall_valueNext;
      case(io_apb_PADDR)
        24'h0000d4 : begin
          if(bus_doWrite)begin
            _zz_565 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000138 : begin
          if(bus_doWrite)begin
            _zz_566 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h00000c : begin
          if(bus_doWrite)begin
            _zz_567 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h00006c : begin
          if(bus_doWrite)begin
            _zz_568 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001b4 : begin
          if(bus_doWrite)begin
            _zz_569 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000108 : begin
          if(bus_doWrite)begin
            _zz_570 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000140 : begin
          if(bus_doWrite)begin
            _zz_571 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h00007c : begin
          if(bus_doWrite)begin
            _zz_572 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001ec : begin
          if(bus_doWrite)begin
            _zz_573 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001bc : begin
          if(bus_doWrite)begin
            _zz_574 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000120 : begin
          if(bus_doWrite)begin
            _zz_575 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000144 : begin
          if(bus_doWrite)begin
            _zz_576 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000130 : begin
          if(bus_doWrite)begin
            _zz_577 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001b0 : begin
          if(bus_doWrite)begin
            _zz_578 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0000d0 : begin
          if(bus_doWrite)begin
            _zz_579 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000054 : begin
          if(bus_doWrite)begin
            _zz_580 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000114 : begin
          if(bus_doWrite)begin
            _zz_581 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000100 : begin
          if(bus_doWrite)begin
            _zz_582 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001a4 : begin
          if(bus_doWrite)begin
            _zz_583 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000154 : begin
          if(bus_doWrite)begin
            _zz_584 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h00002c : begin
          if(bus_doWrite)begin
            _zz_585 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0000e0 : begin
          if(bus_doWrite)begin
            _zz_586 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000118 : begin
          if(bus_doWrite)begin
            _zz_587 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0000c4 : begin
          if(bus_doWrite)begin
            _zz_588 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000098 : begin
          if(bus_doWrite)begin
            _zz_589 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0000fc : begin
          if(bus_doWrite)begin
            _zz_590 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001a8 : begin
          if(bus_doWrite)begin
            _zz_591 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000150 : begin
          if(bus_doWrite)begin
            _zz_592 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001c0 : begin
          if(bus_doWrite)begin
            _zz_593 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000060 : begin
          if(bus_doWrite)begin
            _zz_594 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h0001f0 : begin
          if(bus_doWrite)begin
            _zz_595 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000124 : begin
          if(bus_doWrite)begin
            _zz_596 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000048 : begin
          if(bus_doWrite)begin
            _zz_597 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h00018c : begin
          if(bus_doWrite)begin
            _zz_598 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h000160 : begin
          if(bus_doWrite)begin
            _zz_599 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h200000 : begin
          if(bus_doWrite)begin
            _zz_600 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h002004 : begin
          if(bus_doWrite)begin
            _zz_601 <= _zz_709[0];
            _zz_615 <= _zz_710[0];
            _zz_622 <= _zz_711[0];
            _zz_624 <= _zz_712[0];
            _zz_625 <= _zz_713[0];
            _zz_626 <= _zz_714[0];
          end
        end
        24'h002008 : begin
          if(bus_doWrite)begin
            _zz_602 <= _zz_715[0];
            _zz_606 <= _zz_716[0];
            _zz_607 <= _zz_717[0];
            _zz_611 <= _zz_718[0];
            _zz_612 <= _zz_719[0];
            _zz_613 <= _zz_720[0];
            _zz_617 <= _zz_721[0];
            _zz_618 <= _zz_722[0];
            _zz_620 <= _zz_723[0];
            _zz_623 <= _zz_724[0];
            _zz_628 <= _zz_725[0];
            _zz_632 <= _zz_726[0];
            _zz_635 <= _zz_727[0];
          end
        end
        24'h002000 : begin
          if(bus_doWrite)begin
            _zz_603 <= _zz_728[0];
            _zz_604 <= _zz_729[0];
            _zz_608 <= _zz_730[0];
            _zz_616 <= _zz_731[0];
            _zz_621 <= _zz_732[0];
            _zz_630 <= _zz_733[0];
            _zz_633 <= _zz_734[0];
          end
        end
        24'h00200c : begin
          if(bus_doWrite)begin
            _zz_605 <= _zz_735[0];
            _zz_609 <= _zz_736[0];
            _zz_610 <= _zz_737[0];
            _zz_614 <= _zz_738[0];
            _zz_619 <= _zz_739[0];
            _zz_627 <= _zz_740[0];
            _zz_629 <= _zz_741[0];
            _zz_631 <= _zz_742[0];
            _zz_634 <= _zz_743[0];
          end
        end
        24'h201000 : begin
          if(bus_doWrite)begin
            _zz_636 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h002084 : begin
          if(bus_doWrite)begin
            _zz_637 <= _zz_744[0];
            _zz_651 <= _zz_745[0];
            _zz_658 <= _zz_746[0];
            _zz_660 <= _zz_747[0];
            _zz_661 <= _zz_748[0];
            _zz_662 <= _zz_749[0];
          end
        end
        24'h002088 : begin
          if(bus_doWrite)begin
            _zz_638 <= _zz_750[0];
            _zz_642 <= _zz_751[0];
            _zz_643 <= _zz_752[0];
            _zz_647 <= _zz_753[0];
            _zz_648 <= _zz_754[0];
            _zz_649 <= _zz_755[0];
            _zz_653 <= _zz_756[0];
            _zz_654 <= _zz_757[0];
            _zz_656 <= _zz_758[0];
            _zz_659 <= _zz_759[0];
            _zz_664 <= _zz_760[0];
            _zz_668 <= _zz_761[0];
            _zz_671 <= _zz_762[0];
          end
        end
        24'h002080 : begin
          if(bus_doWrite)begin
            _zz_639 <= _zz_763[0];
            _zz_640 <= _zz_764[0];
            _zz_644 <= _zz_765[0];
            _zz_652 <= _zz_766[0];
            _zz_657 <= _zz_767[0];
            _zz_666 <= _zz_768[0];
            _zz_669 <= _zz_769[0];
          end
        end
        24'h00208c : begin
          if(bus_doWrite)begin
            _zz_641 <= _zz_770[0];
            _zz_645 <= _zz_771[0];
            _zz_646 <= _zz_772[0];
            _zz_650 <= _zz_773[0];
            _zz_655 <= _zz_774[0];
            _zz_663 <= _zz_775[0];
            _zz_665 <= _zz_776[0];
            _zz_667 <= _zz_777[0];
            _zz_670 <= _zz_778[0];
          end
        end
        24'h202000 : begin
          if(bus_doWrite)begin
            _zz_672 <= io_apb_PWDATA[1 : 0];
          end
        end
        24'h002104 : begin
          if(bus_doWrite)begin
            _zz_673 <= _zz_779[0];
            _zz_687 <= _zz_780[0];
            _zz_694 <= _zz_781[0];
            _zz_696 <= _zz_782[0];
            _zz_697 <= _zz_783[0];
            _zz_698 <= _zz_784[0];
          end
        end
        24'h002108 : begin
          if(bus_doWrite)begin
            _zz_674 <= _zz_785[0];
            _zz_678 <= _zz_786[0];
            _zz_679 <= _zz_787[0];
            _zz_683 <= _zz_788[0];
            _zz_684 <= _zz_789[0];
            _zz_685 <= _zz_790[0];
            _zz_689 <= _zz_791[0];
            _zz_690 <= _zz_792[0];
            _zz_692 <= _zz_793[0];
            _zz_695 <= _zz_794[0];
            _zz_700 <= _zz_795[0];
            _zz_704 <= _zz_796[0];
            _zz_707 <= _zz_797[0];
          end
        end
        24'h002100 : begin
          if(bus_doWrite)begin
            _zz_675 <= _zz_798[0];
            _zz_676 <= _zz_799[0];
            _zz_680 <= _zz_800[0];
            _zz_688 <= _zz_801[0];
            _zz_693 <= _zz_802[0];
            _zz_702 <= _zz_803[0];
            _zz_705 <= _zz_804[0];
          end
        end
        24'h00210c : begin
          if(bus_doWrite)begin
            _zz_677 <= _zz_805[0];
            _zz_681 <= _zz_806[0];
            _zz_682 <= _zz_807[0];
            _zz_686 <= _zz_808[0];
            _zz_691 <= _zz_809[0];
            _zz_699 <= _zz_810[0];
            _zz_701 <= _zz_811[0];
            _zz_703 <= _zz_812[0];
            _zz_706 <= _zz_813[0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @ (posedge clk) begin
    targets_0_bestRequest_priority <= (_zz_138 ? _zz_136 : _zz_115);
    targets_0_bestRequest_id <= (_zz_138 ? (_zz_135 ? (_zz_129 ? (_zz_117 ? _zz_814 : _zz_815) : (_zz_120 ? _zz_816 : _zz_817)) : (_zz_132 ? (_zz_123 ? _zz_818 : _zz_819) : (_zz_126 ? _zz_820 : _zz_821))) : (_zz_114 ? (_zz_84 ? targets_0_requests_32_id : targets_0_requests_33_id) : (_zz_87 ? targets_0_requests_34_id : targets_0_requests_35_id)));
    targets_0_bestRequest_valid <= (_zz_138 ? _zz_137 : _zz_116);
    _zz_348 <= (_zz_347 ? _zz_346 : _zz_326);
    _zz_349 <= (_zz_347 ? (_zz_345 ? (_zz_339 ? (_zz_327 ? _zz_822 : _zz_823) : (_zz_330 ? _zz_824 : _zz_825)) : (_zz_342 ? (_zz_333 ? _zz_826 : _zz_827) : (_zz_336 ? _zz_828 : _zz_829))) : (_zz_325 ? (_zz_295 ? 7'h6f : 7'h70) : (_zz_298 ? 7'h7b : 7'h7c)));
    _zz_561 <= (_zz_560 ? _zz_559 : _zz_539);
    _zz_562 <= (_zz_560 ? (_zz_558 ? (_zz_552 ? (_zz_540 ? _zz_862 : _zz_863) : (_zz_543 ? _zz_864 : _zz_865)) : (_zz_555 ? (_zz_546 ? _zz_866 : _zz_867) : (_zz_549 ? _zz_868 : _zz_869))) : (_zz_538 ? (_zz_508 ? 7'h6f : 7'h70) : (_zz_511 ? 7'h7b : 7'h7c)));
  end


endmodule
