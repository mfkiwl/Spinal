// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : unnamed
// Git hash  : adf552d8f500e7419fff395b7049228e4bc5de26



module unnamed (
  input      [10:0]   input_1,
  output     [0:0]    output_0,
  output     [1:0]    output_1,
  output     [1:0]    output_2,
  output     [2:0]    output_3,
  output     [2:0]    output_4,
  output     [2:0]    output_5,
  output     [2:0]    output_6,
  output     [3:0]    output_7,
  output     [3:0]    output_8,
  output     [3:0]    output_9,
  output     [3:0]    output_10
);
  reg        [0:0]    _zz_75;
  reg        [1:0]    _zz_76;
  reg        [1:0]    _zz_77;
  reg        [2:0]    _zz_78;
  reg        [2:0]    _zz_79;
  reg        [2:0]    _zz_80;
  reg        [2:0]    _zz_81;
  reg        [2:0]    _zz_82;
  reg        [2:0]    _zz_83;
  reg        [2:0]    _zz_84;
  reg        [2:0]    _zz_85;
  reg        [2:0]    _zz_86;
  reg        [3:0]    _zz_87;
  reg        [3:0]    _zz_88;
  reg        [3:0]    _zz_89;
  reg        [3:0]    _zz_90;
  reg        [3:0]    _zz_91;
  reg        [3:0]    _zz_92;
  reg        [3:0]    _zz_93;
  reg        [3:0]    _zz_94;
  reg        [3:0]    _zz_95;
  reg        [3:0]    _zz_96;
  reg        [3:0]    _zz_97;
  reg        [3:0]    _zz_98;
  reg        [3:0]    _zz_99;
  reg        [3:0]    _zz_100;
  wire       [0:0]    _zz_101;
  wire       [2:0]    _zz_102;
  wire       [1:0]    _zz_103;
  wire       [2:0]    _zz_104;
  wire       [2:0]    _zz_105;
  wire       [0:0]    _zz_106;
  wire       [2:0]    _zz_107;
  wire       [3:0]    _zz_108;
  wire       [1:0]    _zz_109;
  wire       [2:0]    _zz_110;
  wire       [3:0]    _zz_111;
  wire       [3:0]    _zz_112;
  wire       [3:0]    _zz_113;
  wire       [0:0]    _zz_114;
  wire       [2:0]    _zz_115;
  wire       [3:0]    _zz_116;
  wire       [3:0]    _zz_117;
  wire       [1:0]    _zz_118;
  wire       [2:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [1:0]    _zz_121;
  wire       [2:0]    _zz_122;
  wire       [2:0]    _zz_123;
  wire       [2:0]    _zz_124;
  wire       [2:0]    _zz_125;
  wire       [2:0]    _zz_126;
  wire       [2:0]    _zz_127;
  wire       [2:0]    _zz_128;
  wire       [2:0]    _zz_129;
  wire       [2:0]    _zz_130;
  wire       [2:0]    _zz_131;
  wire       [2:0]    _zz_132;
  wire       [2:0]    _zz_133;
  wire       [2:0]    _zz_134;
  wire       [2:0]    _zz_135;
  wire       [2:0]    _zz_136;
  wire       [2:0]    _zz_137;
  wire       [2:0]    _zz_138;
  wire       [2:0]    _zz_139;
  wire                _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire       [2:0]    _zz_11;
  wire       [2:0]    _zz_12;
  wire       [2:0]    _zz_13;
  wire       [2:0]    _zz_14;
  wire       [2:0]    _zz_15;
  wire       [2:0]    _zz_16;
  wire       [2:0]    _zz_17;
  wire       [2:0]    _zz_18;
  wire       [2:0]    _zz_19;
  wire       [2:0]    _zz_20;
  wire       [2:0]    _zz_21;
  wire       [2:0]    _zz_22;
  wire       [2:0]    _zz_23;
  wire       [2:0]    _zz_24;
  wire       [2:0]    _zz_25;
  wire       [2:0]    _zz_26;
  wire       [2:0]    _zz_27;
  wire       [2:0]    _zz_28;
  wire       [2:0]    _zz_29;
  wire       [2:0]    _zz_30;
  wire       [2:0]    _zz_31;
  wire       [2:0]    _zz_32;
  wire       [2:0]    _zz_33;
  wire       [2:0]    _zz_34;
  wire       [2:0]    _zz_35;
  wire       [2:0]    _zz_36;
  wire       [2:0]    _zz_37;
  wire       [2:0]    _zz_38;
  wire       [2:0]    _zz_39;
  wire       [2:0]    _zz_40;
  wire       [2:0]    _zz_41;
  wire       [2:0]    _zz_42;
  wire       [3:0]    _zz_43;
  wire       [3:0]    _zz_44;
  wire       [3:0]    _zz_45;
  wire       [3:0]    _zz_46;
  wire       [3:0]    _zz_47;
  wire       [3:0]    _zz_48;
  wire       [3:0]    _zz_49;
  wire       [3:0]    _zz_50;
  wire       [3:0]    _zz_51;
  wire       [3:0]    _zz_52;
  wire       [3:0]    _zz_53;
  wire       [3:0]    _zz_54;
  wire       [3:0]    _zz_55;
  wire       [3:0]    _zz_56;
  wire       [3:0]    _zz_57;
  wire       [3:0]    _zz_58;
  wire       [3:0]    _zz_59;
  wire       [3:0]    _zz_60;
  wire       [3:0]    _zz_61;
  wire       [3:0]    _zz_62;
  wire       [3:0]    _zz_63;
  wire       [3:0]    _zz_64;
  wire       [3:0]    _zz_65;
  wire       [3:0]    _zz_66;
  wire       [3:0]    _zz_67;
  wire       [3:0]    _zz_68;
  wire       [3:0]    _zz_69;
  wire       [3:0]    _zz_70;
  wire       [3:0]    _zz_71;
  wire       [3:0]    _zz_72;
  wire       [3:0]    _zz_73;
  wire       [3:0]    _zz_74;

  assign _zz_101 = _zz_4;
  assign _zz_102 = {2'd0, _zz_101};
  assign _zz_103 = {_zz_5,_zz_4};
  assign _zz_104 = {1'd0, _zz_103};
  assign _zz_105 = (_zz_84 + _zz_85);
  assign _zz_106 = _zz_7;
  assign _zz_107 = {2'd0, _zz_106};
  assign _zz_108 = (_zz_87 + _zz_88);
  assign _zz_109 = {_zz_8,_zz_7};
  assign _zz_110 = {1'd0, _zz_109};
  assign _zz_111 = (_zz_90 + _zz_91);
  assign _zz_112 = (_zz_93 + _zz_94);
  assign _zz_113 = (_zz_95 + _zz_96);
  assign _zz_114 = _zz_10;
  assign _zz_115 = {2'd0, _zz_114};
  assign _zz_116 = (_zz_97 + _zz_98);
  assign _zz_117 = (_zz_99 + _zz_100);
  assign _zz_118 = {input_1[10],_zz_10};
  assign _zz_119 = {1'd0, _zz_118};
  assign _zz_120 = _zz_1;
  assign _zz_121 = {_zz_2,_zz_1};
  assign _zz_122 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_123 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_124 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_125 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_126 = {_zz_6,{_zz_5,_zz_4}};
  assign _zz_127 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_128 = {_zz_6,{_zz_5,_zz_4}};
  assign _zz_129 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_130 = {_zz_6,{_zz_5,_zz_4}};
  assign _zz_131 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_132 = {_zz_6,{_zz_5,_zz_4}};
  assign _zz_133 = {_zz_9,{_zz_8,_zz_7}};
  assign _zz_134 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_135 = {_zz_6,{_zz_5,_zz_4}};
  assign _zz_136 = {_zz_9,{_zz_8,_zz_7}};
  assign _zz_137 = {_zz_3,{_zz_2,_zz_1}};
  assign _zz_138 = {_zz_6,{_zz_5,_zz_4}};
  assign _zz_139 = {_zz_9,{_zz_8,_zz_7}};
  always @(*) begin
    case(_zz_120)
      1'b0 : begin
        _zz_75 = 1'b0;
      end
      default : begin
        _zz_75 = 1'b1;
      end
    endcase
  end

  always @(*) begin
    case(_zz_121)
      2'b00 : begin
        _zz_76 = 2'b00;
      end
      2'b01 : begin
        _zz_76 = 2'b01;
      end
      2'b10 : begin
        _zz_76 = 2'b01;
      end
      default : begin
        _zz_76 = 2'b10;
      end
    endcase
  end

  always @(*) begin
    case(_zz_122)
      3'b000 : begin
        _zz_77 = 2'b00;
      end
      3'b001 : begin
        _zz_77 = 2'b01;
      end
      3'b010 : begin
        _zz_77 = 2'b01;
      end
      3'b011 : begin
        _zz_77 = 2'b10;
      end
      3'b100 : begin
        _zz_77 = 2'b01;
      end
      3'b101 : begin
        _zz_77 = 2'b10;
      end
      3'b110 : begin
        _zz_77 = 2'b10;
      end
      default : begin
        _zz_77 = 2'b11;
      end
    endcase
  end

  always @(*) begin
    case(_zz_123)
      3'b000 : begin
        _zz_78 = _zz_11;
      end
      3'b001 : begin
        _zz_78 = _zz_12;
      end
      3'b010 : begin
        _zz_78 = _zz_13;
      end
      3'b011 : begin
        _zz_78 = _zz_14;
      end
      3'b100 : begin
        _zz_78 = _zz_15;
      end
      3'b101 : begin
        _zz_78 = _zz_16;
      end
      3'b110 : begin
        _zz_78 = _zz_17;
      end
      default : begin
        _zz_78 = _zz_18;
      end
    endcase
  end

  always @(*) begin
    case(_zz_102)
      3'b000 : begin
        _zz_79 = _zz_11;
      end
      3'b001 : begin
        _zz_79 = _zz_12;
      end
      3'b010 : begin
        _zz_79 = _zz_13;
      end
      3'b011 : begin
        _zz_79 = _zz_14;
      end
      3'b100 : begin
        _zz_79 = _zz_15;
      end
      3'b101 : begin
        _zz_79 = _zz_16;
      end
      3'b110 : begin
        _zz_79 = _zz_17;
      end
      default : begin
        _zz_79 = _zz_18;
      end
    endcase
  end

  always @(*) begin
    case(_zz_124)
      3'b000 : begin
        _zz_80 = _zz_19;
      end
      3'b001 : begin
        _zz_80 = _zz_20;
      end
      3'b010 : begin
        _zz_80 = _zz_21;
      end
      3'b011 : begin
        _zz_80 = _zz_22;
      end
      3'b100 : begin
        _zz_80 = _zz_23;
      end
      3'b101 : begin
        _zz_80 = _zz_24;
      end
      3'b110 : begin
        _zz_80 = _zz_25;
      end
      default : begin
        _zz_80 = _zz_26;
      end
    endcase
  end

  always @(*) begin
    case(_zz_104)
      3'b000 : begin
        _zz_81 = _zz_19;
      end
      3'b001 : begin
        _zz_81 = _zz_20;
      end
      3'b010 : begin
        _zz_81 = _zz_21;
      end
      3'b011 : begin
        _zz_81 = _zz_22;
      end
      3'b100 : begin
        _zz_81 = _zz_23;
      end
      3'b101 : begin
        _zz_81 = _zz_24;
      end
      3'b110 : begin
        _zz_81 = _zz_25;
      end
      default : begin
        _zz_81 = _zz_26;
      end
    endcase
  end

  always @(*) begin
    case(_zz_125)
      3'b000 : begin
        _zz_82 = _zz_27;
      end
      3'b001 : begin
        _zz_82 = _zz_28;
      end
      3'b010 : begin
        _zz_82 = _zz_29;
      end
      3'b011 : begin
        _zz_82 = _zz_30;
      end
      3'b100 : begin
        _zz_82 = _zz_31;
      end
      3'b101 : begin
        _zz_82 = _zz_32;
      end
      3'b110 : begin
        _zz_82 = _zz_33;
      end
      default : begin
        _zz_82 = _zz_34;
      end
    endcase
  end

  always @(*) begin
    case(_zz_126)
      3'b000 : begin
        _zz_83 = _zz_27;
      end
      3'b001 : begin
        _zz_83 = _zz_28;
      end
      3'b010 : begin
        _zz_83 = _zz_29;
      end
      3'b011 : begin
        _zz_83 = _zz_30;
      end
      3'b100 : begin
        _zz_83 = _zz_31;
      end
      3'b101 : begin
        _zz_83 = _zz_32;
      end
      3'b110 : begin
        _zz_83 = _zz_33;
      end
      default : begin
        _zz_83 = _zz_34;
      end
    endcase
  end

  always @(*) begin
    case(_zz_127)
      3'b000 : begin
        _zz_84 = _zz_35;
      end
      3'b001 : begin
        _zz_84 = _zz_36;
      end
      3'b010 : begin
        _zz_84 = _zz_37;
      end
      3'b011 : begin
        _zz_84 = _zz_38;
      end
      3'b100 : begin
        _zz_84 = _zz_39;
      end
      3'b101 : begin
        _zz_84 = _zz_40;
      end
      3'b110 : begin
        _zz_84 = _zz_41;
      end
      default : begin
        _zz_84 = _zz_42;
      end
    endcase
  end

  always @(*) begin
    case(_zz_128)
      3'b000 : begin
        _zz_85 = _zz_35;
      end
      3'b001 : begin
        _zz_85 = _zz_36;
      end
      3'b010 : begin
        _zz_85 = _zz_37;
      end
      3'b011 : begin
        _zz_85 = _zz_38;
      end
      3'b100 : begin
        _zz_85 = _zz_39;
      end
      3'b101 : begin
        _zz_85 = _zz_40;
      end
      3'b110 : begin
        _zz_85 = _zz_41;
      end
      default : begin
        _zz_85 = _zz_42;
      end
    endcase
  end

  always @(*) begin
    case(_zz_107)
      3'b000 : begin
        _zz_86 = _zz_35;
      end
      3'b001 : begin
        _zz_86 = _zz_36;
      end
      3'b010 : begin
        _zz_86 = _zz_37;
      end
      3'b011 : begin
        _zz_86 = _zz_38;
      end
      3'b100 : begin
        _zz_86 = _zz_39;
      end
      3'b101 : begin
        _zz_86 = _zz_40;
      end
      3'b110 : begin
        _zz_86 = _zz_41;
      end
      default : begin
        _zz_86 = _zz_42;
      end
    endcase
  end

  always @(*) begin
    case(_zz_129)
      3'b000 : begin
        _zz_87 = _zz_43;
      end
      3'b001 : begin
        _zz_87 = _zz_44;
      end
      3'b010 : begin
        _zz_87 = _zz_45;
      end
      3'b011 : begin
        _zz_87 = _zz_46;
      end
      3'b100 : begin
        _zz_87 = _zz_47;
      end
      3'b101 : begin
        _zz_87 = _zz_48;
      end
      3'b110 : begin
        _zz_87 = _zz_49;
      end
      default : begin
        _zz_87 = _zz_50;
      end
    endcase
  end

  always @(*) begin
    case(_zz_130)
      3'b000 : begin
        _zz_88 = _zz_43;
      end
      3'b001 : begin
        _zz_88 = _zz_44;
      end
      3'b010 : begin
        _zz_88 = _zz_45;
      end
      3'b011 : begin
        _zz_88 = _zz_46;
      end
      3'b100 : begin
        _zz_88 = _zz_47;
      end
      3'b101 : begin
        _zz_88 = _zz_48;
      end
      3'b110 : begin
        _zz_88 = _zz_49;
      end
      default : begin
        _zz_88 = _zz_50;
      end
    endcase
  end

  always @(*) begin
    case(_zz_110)
      3'b000 : begin
        _zz_89 = _zz_43;
      end
      3'b001 : begin
        _zz_89 = _zz_44;
      end
      3'b010 : begin
        _zz_89 = _zz_45;
      end
      3'b011 : begin
        _zz_89 = _zz_46;
      end
      3'b100 : begin
        _zz_89 = _zz_47;
      end
      3'b101 : begin
        _zz_89 = _zz_48;
      end
      3'b110 : begin
        _zz_89 = _zz_49;
      end
      default : begin
        _zz_89 = _zz_50;
      end
    endcase
  end

  always @(*) begin
    case(_zz_131)
      3'b000 : begin
        _zz_90 = _zz_51;
      end
      3'b001 : begin
        _zz_90 = _zz_52;
      end
      3'b010 : begin
        _zz_90 = _zz_53;
      end
      3'b011 : begin
        _zz_90 = _zz_54;
      end
      3'b100 : begin
        _zz_90 = _zz_55;
      end
      3'b101 : begin
        _zz_90 = _zz_56;
      end
      3'b110 : begin
        _zz_90 = _zz_57;
      end
      default : begin
        _zz_90 = _zz_58;
      end
    endcase
  end

  always @(*) begin
    case(_zz_132)
      3'b000 : begin
        _zz_91 = _zz_51;
      end
      3'b001 : begin
        _zz_91 = _zz_52;
      end
      3'b010 : begin
        _zz_91 = _zz_53;
      end
      3'b011 : begin
        _zz_91 = _zz_54;
      end
      3'b100 : begin
        _zz_91 = _zz_55;
      end
      3'b101 : begin
        _zz_91 = _zz_56;
      end
      3'b110 : begin
        _zz_91 = _zz_57;
      end
      default : begin
        _zz_91 = _zz_58;
      end
    endcase
  end

  always @(*) begin
    case(_zz_133)
      3'b000 : begin
        _zz_92 = _zz_51;
      end
      3'b001 : begin
        _zz_92 = _zz_52;
      end
      3'b010 : begin
        _zz_92 = _zz_53;
      end
      3'b011 : begin
        _zz_92 = _zz_54;
      end
      3'b100 : begin
        _zz_92 = _zz_55;
      end
      3'b101 : begin
        _zz_92 = _zz_56;
      end
      3'b110 : begin
        _zz_92 = _zz_57;
      end
      default : begin
        _zz_92 = _zz_58;
      end
    endcase
  end

  always @(*) begin
    case(_zz_134)
      3'b000 : begin
        _zz_93 = _zz_59;
      end
      3'b001 : begin
        _zz_93 = _zz_60;
      end
      3'b010 : begin
        _zz_93 = _zz_61;
      end
      3'b011 : begin
        _zz_93 = _zz_62;
      end
      3'b100 : begin
        _zz_93 = _zz_63;
      end
      3'b101 : begin
        _zz_93 = _zz_64;
      end
      3'b110 : begin
        _zz_93 = _zz_65;
      end
      default : begin
        _zz_93 = _zz_66;
      end
    endcase
  end

  always @(*) begin
    case(_zz_135)
      3'b000 : begin
        _zz_94 = _zz_59;
      end
      3'b001 : begin
        _zz_94 = _zz_60;
      end
      3'b010 : begin
        _zz_94 = _zz_61;
      end
      3'b011 : begin
        _zz_94 = _zz_62;
      end
      3'b100 : begin
        _zz_94 = _zz_63;
      end
      3'b101 : begin
        _zz_94 = _zz_64;
      end
      3'b110 : begin
        _zz_94 = _zz_65;
      end
      default : begin
        _zz_94 = _zz_66;
      end
    endcase
  end

  always @(*) begin
    case(_zz_136)
      3'b000 : begin
        _zz_95 = _zz_59;
      end
      3'b001 : begin
        _zz_95 = _zz_60;
      end
      3'b010 : begin
        _zz_95 = _zz_61;
      end
      3'b011 : begin
        _zz_95 = _zz_62;
      end
      3'b100 : begin
        _zz_95 = _zz_63;
      end
      3'b101 : begin
        _zz_95 = _zz_64;
      end
      3'b110 : begin
        _zz_95 = _zz_65;
      end
      default : begin
        _zz_95 = _zz_66;
      end
    endcase
  end

  always @(*) begin
    case(_zz_115)
      3'b000 : begin
        _zz_96 = _zz_59;
      end
      3'b001 : begin
        _zz_96 = _zz_60;
      end
      3'b010 : begin
        _zz_96 = _zz_61;
      end
      3'b011 : begin
        _zz_96 = _zz_62;
      end
      3'b100 : begin
        _zz_96 = _zz_63;
      end
      3'b101 : begin
        _zz_96 = _zz_64;
      end
      3'b110 : begin
        _zz_96 = _zz_65;
      end
      default : begin
        _zz_96 = _zz_66;
      end
    endcase
  end

  always @(*) begin
    case(_zz_137)
      3'b000 : begin
        _zz_97 = _zz_67;
      end
      3'b001 : begin
        _zz_97 = _zz_68;
      end
      3'b010 : begin
        _zz_97 = _zz_69;
      end
      3'b011 : begin
        _zz_97 = _zz_70;
      end
      3'b100 : begin
        _zz_97 = _zz_71;
      end
      3'b101 : begin
        _zz_97 = _zz_72;
      end
      3'b110 : begin
        _zz_97 = _zz_73;
      end
      default : begin
        _zz_97 = _zz_74;
      end
    endcase
  end

  always @(*) begin
    case(_zz_138)
      3'b000 : begin
        _zz_98 = _zz_67;
      end
      3'b001 : begin
        _zz_98 = _zz_68;
      end
      3'b010 : begin
        _zz_98 = _zz_69;
      end
      3'b011 : begin
        _zz_98 = _zz_70;
      end
      3'b100 : begin
        _zz_98 = _zz_71;
      end
      3'b101 : begin
        _zz_98 = _zz_72;
      end
      3'b110 : begin
        _zz_98 = _zz_73;
      end
      default : begin
        _zz_98 = _zz_74;
      end
    endcase
  end

  always @(*) begin
    case(_zz_139)
      3'b000 : begin
        _zz_99 = _zz_67;
      end
      3'b001 : begin
        _zz_99 = _zz_68;
      end
      3'b010 : begin
        _zz_99 = _zz_69;
      end
      3'b011 : begin
        _zz_99 = _zz_70;
      end
      3'b100 : begin
        _zz_99 = _zz_71;
      end
      3'b101 : begin
        _zz_99 = _zz_72;
      end
      3'b110 : begin
        _zz_99 = _zz_73;
      end
      default : begin
        _zz_99 = _zz_74;
      end
    endcase
  end

  always @(*) begin
    case(_zz_119)
      3'b000 : begin
        _zz_100 = _zz_67;
      end
      3'b001 : begin
        _zz_100 = _zz_68;
      end
      3'b010 : begin
        _zz_100 = _zz_69;
      end
      3'b011 : begin
        _zz_100 = _zz_70;
      end
      3'b100 : begin
        _zz_100 = _zz_71;
      end
      3'b101 : begin
        _zz_100 = _zz_72;
      end
      3'b110 : begin
        _zz_100 = _zz_73;
      end
      default : begin
        _zz_100 = _zz_74;
      end
    endcase
  end

  assign _zz_1 = input_1[0];
  assign _zz_2 = input_1[1];
  assign _zz_3 = input_1[2];
  assign _zz_4 = input_1[3];
  assign _zz_5 = input_1[4];
  assign _zz_6 = input_1[5];
  assign _zz_7 = input_1[6];
  assign _zz_8 = input_1[7];
  assign _zz_9 = input_1[8];
  assign _zz_10 = input_1[9];
  assign output_0 = _zz_75;
  assign output_1 = _zz_76;
  assign output_2 = _zz_77;
  assign _zz_11 = 3'b000;
  assign _zz_12 = 3'b001;
  assign _zz_13 = 3'b001;
  assign _zz_14 = 3'b010;
  assign _zz_15 = 3'b001;
  assign _zz_16 = 3'b010;
  assign _zz_17 = 3'b010;
  assign _zz_18 = 3'b011;
  assign output_3 = (_zz_78 + _zz_79);
  assign _zz_19 = 3'b000;
  assign _zz_20 = 3'b001;
  assign _zz_21 = 3'b001;
  assign _zz_22 = 3'b010;
  assign _zz_23 = 3'b001;
  assign _zz_24 = 3'b010;
  assign _zz_25 = 3'b010;
  assign _zz_26 = 3'b011;
  assign output_4 = (_zz_80 + _zz_81);
  assign _zz_27 = 3'b000;
  assign _zz_28 = 3'b001;
  assign _zz_29 = 3'b001;
  assign _zz_30 = 3'b010;
  assign _zz_31 = 3'b001;
  assign _zz_32 = 3'b010;
  assign _zz_33 = 3'b010;
  assign _zz_34 = 3'b011;
  assign output_5 = (_zz_82 + _zz_83);
  assign _zz_35 = 3'b000;
  assign _zz_36 = 3'b001;
  assign _zz_37 = 3'b001;
  assign _zz_38 = 3'b010;
  assign _zz_39 = 3'b001;
  assign _zz_40 = 3'b010;
  assign _zz_41 = 3'b010;
  assign _zz_42 = 3'b011;
  assign output_6 = (_zz_105 + _zz_86);
  assign _zz_43 = 4'b0000;
  assign _zz_44 = 4'b0001;
  assign _zz_45 = 4'b0001;
  assign _zz_46 = 4'b0010;
  assign _zz_47 = 4'b0001;
  assign _zz_48 = 4'b0010;
  assign _zz_49 = 4'b0010;
  assign _zz_50 = 4'b0011;
  assign output_7 = (_zz_108 + _zz_89);
  assign _zz_51 = 4'b0000;
  assign _zz_52 = 4'b0001;
  assign _zz_53 = 4'b0001;
  assign _zz_54 = 4'b0010;
  assign _zz_55 = 4'b0001;
  assign _zz_56 = 4'b0010;
  assign _zz_57 = 4'b0010;
  assign _zz_58 = 4'b0011;
  assign output_8 = (_zz_111 + _zz_92);
  assign _zz_59 = 4'b0000;
  assign _zz_60 = 4'b0001;
  assign _zz_61 = 4'b0001;
  assign _zz_62 = 4'b0010;
  assign _zz_63 = 4'b0001;
  assign _zz_64 = 4'b0010;
  assign _zz_65 = 4'b0010;
  assign _zz_66 = 4'b0011;
  assign output_9 = (_zz_112 + _zz_113);
  assign _zz_67 = 4'b0000;
  assign _zz_68 = 4'b0001;
  assign _zz_69 = 4'b0001;
  assign _zz_70 = 4'b0010;
  assign _zz_71 = 4'b0001;
  assign _zz_72 = 4'b0010;
  assign _zz_73 = 4'b0010;
  assign _zz_74 = 4'b0011;
  assign output_10 = (_zz_116 + _zz_117);

endmodule
