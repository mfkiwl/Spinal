// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : unnamed
// Git hash  : adf552d8f500e7419fff395b7049228e4bc5de26



module unnamed (
  output     [30:0]   x,
  output     [62:0]   y,
  output     [127:0]  z
);

  assign x = 31'h12345678;
  assign y = 63'h1234567812345678;
  assign z = 128'h12345678123456781234567812345678;

endmodule
