// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : Top
// Git hash  : b4281f24a3a26be78ad92c641c5fdf50f14fa460



module Top (
  input      [31:0]   _zz_1,
  input      [31:0]   _zz_2,
  output     [31:0]   _zz_3
);

  assign _zz_3 = (_zz_1 + _zz_2);

endmodule
